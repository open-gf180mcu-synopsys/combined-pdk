magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3090 1660
<< nmos >>
rect 230 210 290 380
rect 340 210 400 380
rect 690 210 750 380
rect 850 210 910 380
rect 1020 210 1080 380
rect 1130 210 1190 380
rect 1300 210 1360 380
rect 1410 210 1470 380
rect 1580 210 1640 380
rect 1690 210 1750 380
rect 1860 210 1920 380
rect 2210 210 2270 380
rect 2320 210 2380 380
rect 2670 210 2730 380
rect 2840 210 2900 380
<< pmos >>
rect 200 1110 260 1450
rect 370 1110 430 1450
rect 690 1110 750 1450
rect 850 1110 910 1450
rect 1020 1110 1080 1450
rect 1130 1110 1190 1450
rect 1300 1110 1360 1450
rect 1410 1110 1470 1450
rect 1580 1110 1640 1450
rect 1690 1110 1750 1450
rect 1860 1110 1920 1450
rect 2180 1110 2240 1450
rect 2350 1110 2410 1450
rect 2670 1110 2730 1450
rect 2840 1110 2900 1450
<< ndiff >>
rect 120 318 230 380
rect 120 272 152 318
rect 198 272 230 318
rect 120 210 230 272
rect 290 210 340 380
rect 400 318 500 380
rect 400 272 432 318
rect 478 272 500 318
rect 400 210 500 272
rect 590 318 690 380
rect 590 272 612 318
rect 658 272 690 318
rect 590 210 690 272
rect 750 210 850 380
rect 910 318 1020 380
rect 910 272 942 318
rect 988 272 1020 318
rect 910 210 1020 272
rect 1080 210 1130 380
rect 1190 278 1300 380
rect 1190 232 1222 278
rect 1268 232 1300 278
rect 1190 210 1300 232
rect 1360 210 1410 380
rect 1470 318 1580 380
rect 1470 272 1502 318
rect 1548 272 1580 318
rect 1470 210 1580 272
rect 1640 210 1690 380
rect 1750 318 1860 380
rect 1750 272 1782 318
rect 1828 272 1860 318
rect 1750 210 1860 272
rect 1920 318 2020 380
rect 1920 272 1952 318
rect 1998 272 2020 318
rect 1920 210 2020 272
rect 2110 318 2210 380
rect 2110 272 2132 318
rect 2178 272 2210 318
rect 2110 210 2210 272
rect 2270 210 2320 380
rect 2380 318 2480 380
rect 2380 272 2412 318
rect 2458 272 2480 318
rect 2380 210 2480 272
rect 2570 318 2670 380
rect 2570 272 2592 318
rect 2638 272 2670 318
rect 2570 210 2670 272
rect 2730 318 2840 380
rect 2730 272 2762 318
rect 2808 272 2840 318
rect 2730 210 2840 272
rect 2900 318 3000 380
rect 2900 272 2932 318
rect 2978 272 3000 318
rect 2900 210 3000 272
<< pdiff >>
rect 90 1425 200 1450
rect 90 1285 122 1425
rect 168 1285 200 1425
rect 90 1110 200 1285
rect 260 1425 370 1450
rect 260 1285 292 1425
rect 338 1285 370 1425
rect 260 1110 370 1285
rect 430 1425 530 1450
rect 430 1285 462 1425
rect 508 1285 530 1425
rect 430 1110 530 1285
rect 590 1397 690 1450
rect 590 1163 612 1397
rect 658 1163 690 1397
rect 590 1110 690 1163
rect 750 1110 850 1450
rect 910 1397 1020 1450
rect 910 1163 942 1397
rect 988 1163 1020 1397
rect 910 1110 1020 1163
rect 1080 1110 1130 1450
rect 1190 1397 1300 1450
rect 1190 1163 1222 1397
rect 1268 1163 1300 1397
rect 1190 1110 1300 1163
rect 1360 1110 1410 1450
rect 1470 1425 1580 1450
rect 1470 1285 1502 1425
rect 1548 1285 1580 1425
rect 1470 1110 1580 1285
rect 1640 1110 1690 1450
rect 1750 1425 1860 1450
rect 1750 1285 1782 1425
rect 1828 1285 1860 1425
rect 1750 1110 1860 1285
rect 1920 1397 2020 1450
rect 1920 1163 1952 1397
rect 1998 1163 2020 1397
rect 1920 1110 2020 1163
rect 2080 1430 2180 1450
rect 2080 1290 2102 1430
rect 2148 1290 2180 1430
rect 2080 1110 2180 1290
rect 2240 1428 2350 1450
rect 2240 1382 2272 1428
rect 2318 1382 2350 1428
rect 2240 1110 2350 1382
rect 2410 1388 2510 1450
rect 2410 1342 2442 1388
rect 2488 1342 2510 1388
rect 2410 1110 2510 1342
rect 2570 1397 2670 1450
rect 2570 1163 2592 1397
rect 2638 1163 2670 1397
rect 2570 1110 2670 1163
rect 2730 1397 2840 1450
rect 2730 1163 2762 1397
rect 2808 1163 2840 1397
rect 2730 1110 2840 1163
rect 2900 1397 3000 1450
rect 2900 1163 2932 1397
rect 2978 1163 3000 1397
rect 2900 1110 3000 1163
<< ndiffc >>
rect 152 272 198 318
rect 432 272 478 318
rect 612 272 658 318
rect 942 272 988 318
rect 1222 232 1268 278
rect 1502 272 1548 318
rect 1782 272 1828 318
rect 1952 272 1998 318
rect 2132 272 2178 318
rect 2412 272 2458 318
rect 2592 272 2638 318
rect 2762 272 2808 318
rect 2932 272 2978 318
<< pdiffc >>
rect 122 1285 168 1425
rect 292 1285 338 1425
rect 462 1285 508 1425
rect 612 1163 658 1397
rect 942 1163 988 1397
rect 1222 1163 1268 1397
rect 1502 1285 1548 1425
rect 1782 1285 1828 1425
rect 1952 1163 1998 1397
rect 2102 1290 2148 1430
rect 2272 1382 2318 1428
rect 2442 1342 2488 1388
rect 2592 1163 2638 1397
rect 2762 1163 2808 1397
rect 2932 1163 2978 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
rect 980 118 1130 140
rect 980 72 1032 118
rect 1078 72 1130 118
rect 980 50 1130 72
rect 1210 118 1360 140
rect 1210 72 1262 118
rect 1308 72 1360 118
rect 1210 50 1360 72
rect 1440 118 1590 140
rect 1440 72 1492 118
rect 1538 72 1590 118
rect 1440 50 1590 72
rect 1670 118 1820 140
rect 1670 72 1722 118
rect 1768 72 1820 118
rect 1670 50 1820 72
rect 1900 118 2050 140
rect 1900 72 1952 118
rect 1998 72 2050 118
rect 1900 50 2050 72
rect 2130 118 2280 140
rect 2130 72 2182 118
rect 2228 72 2280 118
rect 2130 50 2280 72
rect 2360 118 2510 140
rect 2360 72 2412 118
rect 2458 72 2510 118
rect 2360 50 2510 72
rect 2590 118 2740 140
rect 2590 72 2642 118
rect 2688 72 2740 118
rect 2590 50 2740 72
rect 2820 118 2970 140
rect 2820 72 2872 118
rect 2918 72 2970 118
rect 2820 50 2970 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
rect 980 1588 1130 1610
rect 980 1542 1032 1588
rect 1078 1542 1130 1588
rect 980 1520 1130 1542
rect 1210 1588 1360 1610
rect 1210 1542 1262 1588
rect 1308 1542 1360 1588
rect 1210 1520 1360 1542
rect 1440 1588 1590 1610
rect 1440 1542 1492 1588
rect 1538 1542 1590 1588
rect 1440 1520 1590 1542
rect 1670 1588 1820 1610
rect 1670 1542 1722 1588
rect 1768 1542 1820 1588
rect 1670 1520 1820 1542
rect 1900 1588 2050 1610
rect 1900 1542 1952 1588
rect 1998 1542 2050 1588
rect 1900 1520 2050 1542
rect 2130 1588 2280 1610
rect 2130 1542 2182 1588
rect 2228 1542 2280 1588
rect 2130 1520 2280 1542
rect 2360 1588 2510 1610
rect 2360 1542 2412 1588
rect 2458 1542 2510 1588
rect 2360 1520 2510 1542
rect 2590 1588 2740 1610
rect 2590 1542 2642 1588
rect 2688 1542 2740 1588
rect 2590 1520 2740 1542
rect 2820 1588 2970 1610
rect 2820 1542 2872 1588
rect 2918 1542 2970 1588
rect 2820 1520 2970 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
rect 1032 72 1078 118
rect 1262 72 1308 118
rect 1492 72 1538 118
rect 1722 72 1768 118
rect 1952 72 1998 118
rect 2182 72 2228 118
rect 2412 72 2458 118
rect 2642 72 2688 118
rect 2872 72 2918 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
rect 1032 1542 1078 1588
rect 1262 1542 1308 1588
rect 1492 1542 1538 1588
rect 1722 1542 1768 1588
rect 1952 1542 1998 1588
rect 2182 1542 2228 1588
rect 2412 1542 2458 1588
rect 2642 1542 2688 1588
rect 2872 1542 2918 1588
<< polysilicon >>
rect 200 1450 260 1500
rect 370 1450 430 1500
rect 690 1450 750 1500
rect 850 1450 910 1500
rect 1020 1450 1080 1500
rect 1130 1450 1190 1500
rect 1300 1450 1360 1500
rect 1410 1450 1470 1500
rect 1580 1450 1640 1500
rect 1690 1450 1750 1500
rect 1860 1450 1920 1500
rect 2180 1450 2240 1500
rect 2350 1450 2410 1500
rect 2670 1450 2730 1500
rect 2840 1450 2900 1500
rect 200 930 260 1110
rect 200 903 320 930
rect 200 857 227 903
rect 273 857 320 903
rect 200 830 320 857
rect 200 470 260 830
rect 370 800 430 1110
rect 690 800 750 1110
rect 850 930 910 1110
rect 850 903 950 930
rect 850 857 877 903
rect 923 857 950 903
rect 850 830 950 857
rect 370 773 510 800
rect 370 727 427 773
rect 473 727 510 773
rect 370 700 510 727
rect 690 773 810 800
rect 690 727 737 773
rect 783 727 810 773
rect 690 700 810 727
rect 370 470 430 700
rect 200 430 290 470
rect 230 380 290 430
rect 340 430 430 470
rect 340 380 400 430
rect 690 380 750 700
rect 1020 660 1080 1110
rect 1130 1060 1190 1110
rect 1300 1060 1360 1110
rect 1130 1033 1360 1060
rect 1130 990 1167 1033
rect 1140 987 1167 990
rect 1213 990 1360 1033
rect 1213 987 1240 990
rect 1140 940 1240 987
rect 1410 660 1470 1110
rect 1580 930 1640 1110
rect 1540 903 1640 930
rect 1540 857 1567 903
rect 1613 857 1640 903
rect 1540 830 1640 857
rect 1690 800 1750 1110
rect 1860 930 1920 1110
rect 1860 903 1960 930
rect 1860 857 1887 903
rect 1933 857 1960 903
rect 1860 830 1960 857
rect 1680 773 1780 800
rect 1680 727 1707 773
rect 1753 727 1780 773
rect 1680 700 1780 727
rect 1540 660 1640 670
rect 850 643 1640 660
rect 850 600 1567 643
rect 850 380 910 600
rect 1540 597 1567 600
rect 1613 597 1640 643
rect 1540 570 1640 597
rect 980 513 1080 540
rect 1140 520 1240 540
rect 980 467 1007 513
rect 1053 467 1080 513
rect 980 440 1080 467
rect 1020 380 1080 440
rect 1130 513 1360 520
rect 1130 467 1167 513
rect 1213 467 1360 513
rect 1130 440 1360 467
rect 1130 380 1190 440
rect 1300 380 1360 440
rect 1410 503 1510 530
rect 1410 457 1437 503
rect 1483 457 1510 503
rect 1410 430 1510 457
rect 1410 380 1470 430
rect 1580 380 1640 570
rect 1690 380 1750 700
rect 1860 380 1920 830
rect 2180 530 2240 1110
rect 2350 930 2410 1110
rect 2290 903 2410 930
rect 2290 857 2337 903
rect 2383 857 2410 903
rect 2290 830 2410 857
rect 2100 503 2240 530
rect 2100 457 2137 503
rect 2183 470 2240 503
rect 2350 470 2410 830
rect 2670 670 2730 1110
rect 2840 930 2900 1110
rect 2780 903 2900 930
rect 2780 857 2807 903
rect 2853 857 2900 903
rect 2780 830 2900 857
rect 2610 643 2730 670
rect 2610 597 2657 643
rect 2703 597 2730 643
rect 2610 570 2730 597
rect 2183 457 2270 470
rect 2100 430 2270 457
rect 2210 380 2270 430
rect 2320 430 2410 470
rect 2320 380 2380 430
rect 2670 380 2730 570
rect 2840 380 2900 830
rect 230 160 290 210
rect 340 160 400 210
rect 690 160 750 210
rect 850 160 910 210
rect 1020 160 1080 210
rect 1130 160 1190 210
rect 1300 160 1360 210
rect 1410 160 1470 210
rect 1580 160 1640 210
rect 1690 160 1750 210
rect 1860 160 1920 210
rect 2210 160 2270 210
rect 2320 160 2380 210
rect 2670 160 2730 210
rect 2840 160 2900 210
<< polycontact >>
rect 227 857 273 903
rect 877 857 923 903
rect 427 727 473 773
rect 737 727 783 773
rect 1167 987 1213 1033
rect 1567 857 1613 903
rect 1887 857 1933 903
rect 1707 727 1753 773
rect 1567 597 1613 643
rect 1007 467 1053 513
rect 1167 467 1213 513
rect 1437 457 1483 503
rect 2337 857 2383 903
rect 2137 457 2183 503
rect 2807 857 2853 903
rect 2657 597 2703 643
<< metal1 >>
rect 0 1588 3090 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1032 1588
rect 1078 1542 1262 1588
rect 1308 1542 1492 1588
rect 1538 1542 1722 1588
rect 1768 1542 1952 1588
rect 1998 1542 2182 1588
rect 2228 1542 2412 1588
rect 2458 1542 2642 1588
rect 2688 1542 2872 1588
rect 2918 1542 3090 1588
rect 0 1520 3090 1542
rect 120 1425 170 1450
rect 120 1285 122 1425
rect 168 1285 170 1425
rect 120 1210 170 1285
rect 290 1425 340 1520
rect 290 1285 292 1425
rect 338 1285 340 1425
rect 290 1260 340 1285
rect 460 1425 510 1450
rect 460 1285 462 1425
rect 508 1285 510 1425
rect 460 1210 510 1285
rect 120 1160 510 1210
rect 610 1397 660 1520
rect 610 1163 612 1397
rect 658 1163 660 1397
rect 150 910 200 1160
rect 610 1110 660 1163
rect 940 1397 990 1450
rect 940 1163 942 1397
rect 988 1163 990 1397
rect 940 1060 990 1163
rect 1220 1397 1270 1520
rect 1220 1163 1222 1397
rect 1268 1163 1270 1397
rect 1500 1425 1550 1450
rect 1500 1285 1502 1425
rect 1548 1285 1550 1425
rect 1500 1260 1550 1285
rect 1780 1425 1830 1520
rect 1780 1285 1782 1425
rect 1828 1285 1830 1425
rect 1780 1260 1830 1285
rect 1950 1397 2000 1450
rect 1220 1110 1270 1163
rect 1320 1210 1550 1260
rect 610 1010 990 1060
rect 1140 1033 1240 1040
rect 150 906 300 910
rect 150 854 224 906
rect 276 854 300 906
rect 150 850 300 854
rect 150 520 200 850
rect 610 780 660 1010
rect 1140 987 1167 1033
rect 1213 987 1240 1033
rect 1140 980 1240 987
rect 850 906 1080 910
rect 850 903 1004 906
rect 850 857 877 903
rect 923 857 1004 903
rect 850 854 1004 857
rect 1056 854 1080 906
rect 850 850 1080 854
rect 400 776 660 780
rect 400 724 424 776
rect 476 724 660 776
rect 400 720 660 724
rect 710 776 810 780
rect 710 724 734 776
rect 786 724 810 776
rect 710 720 810 724
rect 420 520 470 530
rect 610 520 660 720
rect 1000 520 1060 850
rect 1160 520 1220 980
rect 1320 760 1370 1210
rect 1950 1163 1952 1397
rect 1998 1163 2000 1397
rect 2100 1430 2150 1450
rect 2100 1290 2102 1430
rect 2148 1310 2150 1430
rect 2270 1428 2320 1520
rect 2270 1382 2272 1428
rect 2318 1382 2320 1428
rect 2270 1360 2320 1382
rect 2440 1388 2490 1450
rect 2440 1342 2442 1388
rect 2488 1342 2490 1388
rect 2440 1310 2490 1342
rect 2148 1290 2490 1310
rect 2100 1260 2490 1290
rect 2590 1397 2640 1450
rect 1670 1036 1770 1040
rect 1670 984 1694 1036
rect 1746 984 1770 1036
rect 1670 980 1770 984
rect 1950 1020 2000 1163
rect 2590 1163 2592 1397
rect 2638 1163 2640 1397
rect 2130 1040 2190 1060
rect 2470 1040 2530 1060
rect 2130 1036 2530 1040
rect 1310 710 1370 760
rect 1430 906 1640 910
rect 1430 854 1564 906
rect 1616 854 1640 906
rect 1430 850 1640 854
rect 150 516 500 520
rect 150 464 424 516
rect 476 464 500 516
rect 610 470 810 520
rect 150 460 500 464
rect 150 318 200 460
rect 420 450 470 460
rect 730 380 810 470
rect 980 513 1080 520
rect 980 467 1007 513
rect 1053 467 1080 513
rect 980 460 1080 467
rect 1140 516 1240 520
rect 1140 464 1164 516
rect 1216 464 1240 516
rect 1140 460 1240 464
rect 1310 390 1360 710
rect 1430 510 1490 850
rect 1690 780 1750 980
rect 1950 970 2060 1020
rect 1860 906 1960 910
rect 1860 854 1884 906
rect 1936 854 1960 906
rect 1860 850 1960 854
rect 2010 780 2060 970
rect 2130 984 2134 1036
rect 2186 984 2474 1036
rect 2526 984 2530 1036
rect 2130 980 2530 984
rect 2130 960 2190 980
rect 2310 906 2410 910
rect 2310 854 2334 906
rect 2386 854 2410 906
rect 2310 850 2410 854
rect 1680 776 1780 780
rect 1680 724 1704 776
rect 1756 724 1780 776
rect 1680 720 1780 724
rect 1950 730 2060 780
rect 1540 646 1640 650
rect 1540 594 1564 646
rect 1616 594 1640 646
rect 1540 590 1640 594
rect 1950 646 2010 730
rect 2470 650 2530 980
rect 2590 910 2640 1163
rect 2760 1397 2810 1520
rect 2760 1163 2762 1397
rect 2808 1163 2810 1397
rect 2760 1110 2810 1163
rect 2930 1397 2980 1450
rect 2930 1163 2932 1397
rect 2978 1163 2980 1397
rect 2930 1050 2980 1163
rect 2930 1036 3030 1050
rect 2930 984 2954 1036
rect 3006 984 3030 1036
rect 2930 980 3030 984
rect 2930 970 3020 980
rect 2590 906 2880 910
rect 2590 854 2804 906
rect 2856 854 2880 906
rect 2590 850 2880 854
rect 1950 594 1954 646
rect 2006 594 2010 646
rect 1950 570 2010 594
rect 2410 646 2730 650
rect 2410 594 2654 646
rect 2706 594 2730 646
rect 2410 590 2730 594
rect 1410 503 1510 510
rect 1410 457 1437 503
rect 1483 457 1510 503
rect 1410 450 1510 457
rect 1310 386 1580 390
rect 150 272 152 318
rect 198 272 200 318
rect 150 210 200 272
rect 430 318 480 380
rect 430 272 432 318
rect 478 272 480 318
rect 430 140 480 272
rect 610 318 660 380
rect 730 330 990 380
rect 1310 340 1504 386
rect 610 272 612 318
rect 658 272 660 318
rect 610 140 660 272
rect 940 318 990 330
rect 940 272 942 318
rect 988 272 990 318
rect 1500 334 1504 340
rect 1556 334 1580 386
rect 1500 330 1580 334
rect 1500 318 1550 330
rect 940 210 990 272
rect 1220 278 1270 300
rect 1220 232 1222 278
rect 1268 232 1270 278
rect 1220 140 1270 232
rect 1500 272 1502 318
rect 1548 272 1550 318
rect 1500 210 1550 272
rect 1780 318 1830 380
rect 1780 272 1782 318
rect 1828 272 1830 318
rect 1780 140 1830 272
rect 1950 318 2000 570
rect 2110 506 2210 510
rect 2110 454 2134 506
rect 2186 454 2210 506
rect 2110 450 2210 454
rect 1950 272 1952 318
rect 1998 272 2000 318
rect 1950 210 2000 272
rect 2130 318 2180 380
rect 2130 272 2132 318
rect 2178 272 2180 318
rect 2130 140 2180 272
rect 2410 318 2460 590
rect 2810 480 2860 850
rect 2410 272 2412 318
rect 2458 272 2460 318
rect 2410 210 2460 272
rect 2590 430 2860 480
rect 2590 318 2640 430
rect 2590 272 2592 318
rect 2638 272 2640 318
rect 2590 210 2640 272
rect 2760 318 2810 380
rect 2760 272 2762 318
rect 2808 272 2810 318
rect 2760 140 2810 272
rect 2930 318 2980 970
rect 2930 272 2932 318
rect 2978 272 2980 318
rect 2930 210 2980 272
rect 0 118 3090 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1032 118
rect 1078 72 1262 118
rect 1308 72 1492 118
rect 1538 72 1722 118
rect 1768 72 1952 118
rect 1998 72 2182 118
rect 2228 72 2412 118
rect 2458 72 2642 118
rect 2688 72 2872 118
rect 2918 72 3090 118
rect 0 0 3090 72
<< via1 >>
rect 224 903 276 906
rect 224 857 227 903
rect 227 857 273 903
rect 273 857 276 903
rect 224 854 276 857
rect 1004 854 1056 906
rect 424 773 476 776
rect 424 727 427 773
rect 427 727 473 773
rect 473 727 476 773
rect 424 724 476 727
rect 734 773 786 776
rect 734 727 737 773
rect 737 727 783 773
rect 783 727 786 773
rect 734 724 786 727
rect 1694 984 1746 1036
rect 1564 903 1616 906
rect 1564 857 1567 903
rect 1567 857 1613 903
rect 1613 857 1616 903
rect 1564 854 1616 857
rect 424 464 476 516
rect 1164 513 1216 516
rect 1164 467 1167 513
rect 1167 467 1213 513
rect 1213 467 1216 513
rect 1164 464 1216 467
rect 1884 903 1936 906
rect 1884 857 1887 903
rect 1887 857 1933 903
rect 1933 857 1936 903
rect 1884 854 1936 857
rect 2134 984 2186 1036
rect 2474 984 2526 1036
rect 2334 903 2386 906
rect 2334 857 2337 903
rect 2337 857 2383 903
rect 2383 857 2386 903
rect 2334 854 2386 857
rect 1704 773 1756 776
rect 1704 727 1707 773
rect 1707 727 1753 773
rect 1753 727 1756 773
rect 1704 724 1756 727
rect 1564 643 1616 646
rect 1564 597 1567 643
rect 1567 597 1613 643
rect 1613 597 1616 643
rect 1564 594 1616 597
rect 2954 984 3006 1036
rect 2804 903 2856 906
rect 2804 857 2807 903
rect 2807 857 2853 903
rect 2853 857 2856 903
rect 2804 854 2856 857
rect 1954 594 2006 646
rect 2654 643 2706 646
rect 2654 597 2657 643
rect 2657 597 2703 643
rect 2703 597 2706 643
rect 2654 594 2706 597
rect 1504 334 1556 386
rect 2134 503 2186 506
rect 2134 457 2137 503
rect 2137 457 2183 503
rect 2183 457 2186 503
rect 2134 454 2186 457
<< metal2 >>
rect 220 1110 2390 1170
rect 220 920 280 1110
rect 1680 1040 1760 1050
rect 2120 1040 2200 1050
rect 1670 1036 2210 1040
rect 1670 984 1694 1036
rect 1746 984 2134 1036
rect 2186 984 2210 1036
rect 1670 980 2210 984
rect 1680 970 1760 980
rect 2120 970 2200 980
rect 2330 920 2390 1110
rect 2450 1036 2550 1050
rect 2940 1040 3020 1050
rect 2450 984 2474 1036
rect 2526 984 2550 1036
rect 2450 970 2550 984
rect 2930 1036 3030 1040
rect 2930 984 2954 1036
rect 3006 984 3030 1036
rect 2930 980 3030 984
rect 2940 970 3020 980
rect 200 906 300 920
rect 200 854 224 906
rect 276 854 300 906
rect 200 840 300 854
rect 980 910 1070 920
rect 1540 910 1640 920
rect 1870 910 1950 920
rect 980 906 1960 910
rect 980 854 1004 906
rect 1056 854 1564 906
rect 1616 854 1884 906
rect 1936 854 1960 906
rect 980 850 1960 854
rect 2310 906 2410 920
rect 2790 910 2870 920
rect 2310 854 2334 906
rect 2386 854 2410 906
rect 980 840 1070 850
rect 1540 840 1640 850
rect 1870 840 1950 850
rect 2310 840 2410 854
rect 2780 906 2880 910
rect 2780 854 2804 906
rect 2856 854 2880 906
rect 2780 850 2880 854
rect 2790 840 2870 850
rect 400 776 500 790
rect 400 724 424 776
rect 476 724 500 776
rect 400 710 500 724
rect 710 776 810 790
rect 1690 780 1770 790
rect 710 724 734 776
rect 786 724 810 776
rect 710 710 810 724
rect 1680 776 1780 780
rect 1680 724 1704 776
rect 1756 724 1780 776
rect 1680 720 1780 724
rect 1690 710 1770 720
rect 1550 650 1630 660
rect 1940 650 2020 660
rect 2640 650 2720 660
rect 1540 646 2040 650
rect 1540 594 1564 646
rect 1616 594 1954 646
rect 2006 594 2040 646
rect 1540 590 2040 594
rect 2570 646 2730 650
rect 2570 594 2654 646
rect 2706 594 2730 646
rect 2570 590 2730 594
rect 1550 580 1630 590
rect 1940 580 2020 590
rect 2640 580 2720 590
rect 400 520 500 530
rect 1150 520 1230 530
rect 400 516 1240 520
rect 400 464 424 516
rect 476 464 1164 516
rect 1216 464 1240 516
rect 400 460 1240 464
rect 2110 506 2210 520
rect 400 450 500 460
rect 1150 450 1230 460
rect 2110 454 2134 506
rect 2186 454 2210 506
rect 2110 440 2210 454
rect 1490 390 1570 400
rect 2110 390 2190 440
rect 1480 386 2190 390
rect 1480 334 1504 386
rect 1556 334 2190 386
rect 1480 330 2190 334
rect 1490 320 1570 330
<< labels >>
rlabel via1 s 734 724 786 776 4 D
port 1 nsew signal input
rlabel via1 s 2954 984 3006 1036 4 Q
port 2 nsew signal output
rlabel via1 s 2804 854 2856 906 4 QN
port 3 nsew signal output
rlabel via1 s 2334 854 2386 906 4 SN
port 4 nsew signal output
rlabel via1 s 1884 854 1936 906 4 CLK
port 5 nsew clock input
rlabel metal1 s 290 1260 340 1660 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 430 0 480 380 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 610 1110 660 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1220 1110 1270 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1780 1260 1830 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2270 1360 2320 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2760 1110 2810 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3090 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 0 660 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1220 0 1270 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1780 0 1830 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2130 0 2180 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2760 0 2810 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3090 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel via1 s 1564 854 1616 906 1 CLK
port 5 nsew clock input
rlabel via1 s 1004 854 1056 906 1 CLK
port 5 nsew clock input
rlabel metal2 s 980 840 1070 920 1 CLK
port 5 nsew clock input
rlabel metal2 s 1540 840 1640 920 1 CLK
port 5 nsew clock input
rlabel metal2 s 1870 840 1950 920 1 CLK
port 5 nsew clock input
rlabel metal2 s 980 850 1960 910 1 CLK
port 5 nsew clock input
rlabel metal1 s 1000 460 1060 910 1 CLK
port 5 nsew clock input
rlabel metal1 s 980 460 1080 520 1 CLK
port 5 nsew clock input
rlabel metal1 s 850 850 1080 910 1 CLK
port 5 nsew clock input
rlabel metal1 s 1430 450 1490 910 1 CLK
port 5 nsew clock input
rlabel metal1 s 1410 450 1510 510 1 CLK
port 5 nsew clock input
rlabel metal1 s 1430 850 1640 910 1 CLK
port 5 nsew clock input
rlabel metal1 s 1860 850 1960 910 1 CLK
port 5 nsew clock input
rlabel metal2 s 710 710 810 790 1 D
port 1 nsew signal input
rlabel metal1 s 710 720 810 780 1 D
port 1 nsew signal input
rlabel metal2 s 2940 970 3020 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 2930 980 3030 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 2930 210 2980 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 2930 970 3020 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 2930 980 3030 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 2790 840 2870 920 1 QN
port 3 nsew signal output
rlabel metal2 s 2780 850 2880 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2590 210 2640 480 1 QN
port 3 nsew signal output
rlabel metal1 s 2590 850 2640 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 2590 430 2860 480 1 QN
port 3 nsew signal output
rlabel metal1 s 2810 430 2860 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2590 850 2880 910 1 QN
port 3 nsew signal output
rlabel via1 s 1164 464 1216 516 1 SN
port 4 nsew signal output
rlabel via1 s 424 464 476 516 1 SN
port 4 nsew signal output
rlabel via1 s 224 854 276 906 1 SN
port 4 nsew signal output
rlabel metal2 s 400 450 500 530 1 SN
port 4 nsew signal output
rlabel metal2 s 1150 450 1230 530 1 SN
port 4 nsew signal output
rlabel metal2 s 400 460 1240 520 1 SN
port 4 nsew signal output
rlabel metal2 s 220 840 280 1170 1 SN
port 4 nsew signal output
rlabel metal2 s 200 840 300 920 1 SN
port 4 nsew signal output
rlabel metal2 s 2330 840 2390 1170 1 SN
port 4 nsew signal output
rlabel metal2 s 220 1110 2390 1170 1 SN
port 4 nsew signal output
rlabel metal2 s 2310 840 2410 920 1 SN
port 4 nsew signal output
rlabel metal1 s 120 1160 170 1450 1 SN
port 4 nsew signal output
rlabel metal1 s 150 210 200 1210 1 SN
port 4 nsew signal output
rlabel metal1 s 150 850 300 910 1 SN
port 4 nsew signal output
rlabel metal1 s 120 1160 510 1210 1 SN
port 4 nsew signal output
rlabel metal1 s 420 450 470 530 1 SN
port 4 nsew signal output
rlabel metal1 s 150 460 500 520 1 SN
port 4 nsew signal output
rlabel metal1 s 460 1160 510 1450 1 SN
port 4 nsew signal output
rlabel metal1 s 1160 460 1220 1040 1 SN
port 4 nsew signal output
rlabel metal1 s 1140 460 1240 520 1 SN
port 4 nsew signal output
rlabel metal1 s 1140 980 1240 1040 1 SN
port 4 nsew signal output
rlabel metal1 s 2310 850 2410 910 1 SN
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3090 1660
string GDS_END 289962
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 266966
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
