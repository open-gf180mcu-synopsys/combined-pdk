magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 820 1270
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
rect 570 210 630 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 570 720 630 1060
<< ndiff >>
rect 120 278 220 380
rect 120 232 142 278
rect 188 232 220 278
rect 120 210 220 232
rect 280 210 330 380
rect 390 318 570 380
rect 390 272 457 318
rect 503 272 570 318
rect 390 210 570 272
rect 630 278 730 380
rect 630 232 662 278
rect 708 232 730 278
rect 630 210 730 232
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 360 1060
rect 250 773 282 1007
rect 328 773 360 1007
rect 250 720 360 773
rect 420 1007 570 1060
rect 420 773 472 1007
rect 518 773 570 1007
rect 420 720 570 773
rect 630 1013 730 1060
rect 630 967 662 1013
rect 708 967 730 1013
rect 630 720 730 967
<< ndiffc >>
rect 142 232 188 278
rect 457 272 503 318
rect 662 232 708 278
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 472 773 518 1007
rect 662 967 708 1013
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 570 1060 630 1110
rect 190 540 250 720
rect 360 670 420 720
rect 360 643 490 670
rect 360 630 417 643
rect 110 513 250 540
rect 110 467 147 513
rect 193 480 250 513
rect 330 597 417 630
rect 463 597 490 643
rect 330 570 490 597
rect 193 467 280 480
rect 110 440 280 467
rect 220 380 280 440
rect 330 380 390 570
rect 570 540 630 720
rect 530 513 630 540
rect 530 467 557 513
rect 603 467 630 513
rect 530 440 630 467
rect 570 380 630 440
rect 220 160 280 210
rect 330 160 390 210
rect 570 160 630 210
<< polycontact >>
rect 147 467 193 513
rect 417 597 463 643
rect 557 467 603 513
<< metal1 >>
rect 0 1198 820 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 820 1198
rect 0 1130 820 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 520 330 773
rect 450 1007 540 1130
rect 450 773 472 1007
rect 518 773 540 1007
rect 450 720 540 773
rect 660 1013 710 1060
rect 660 967 662 1013
rect 708 967 710 1013
rect 660 790 710 967
rect 660 780 740 790
rect 660 776 760 780
rect 660 724 684 776
rect 736 724 760 776
rect 660 720 760 724
rect 660 710 740 720
rect 390 646 490 650
rect 390 594 414 646
rect 466 594 490 646
rect 390 590 490 594
rect 550 520 610 540
rect 120 516 220 520
rect 120 464 144 516
rect 196 464 220 516
rect 120 460 220 464
rect 280 513 610 520
rect 280 467 557 513
rect 603 467 610 513
rect 280 460 610 467
rect 280 360 330 460
rect 550 440 610 460
rect 140 310 330 360
rect 420 318 540 380
rect 140 278 190 310
rect 140 232 142 278
rect 188 232 190 278
rect 140 210 190 232
rect 420 272 457 318
rect 503 272 540 318
rect 420 140 540 272
rect 660 278 710 710
rect 660 232 662 278
rect 708 232 710 278
rect 660 210 710 232
rect 0 118 820 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 820 118
rect 0 0 820 72
<< via1 >>
rect 684 724 736 776
rect 414 643 466 646
rect 414 597 417 643
rect 417 597 463 643
rect 463 597 466 643
rect 414 594 466 597
rect 144 513 196 516
rect 144 467 147 513
rect 147 467 193 513
rect 193 467 196 513
rect 144 464 196 467
<< metal2 >>
rect 660 776 760 790
rect 660 724 684 776
rect 736 724 760 776
rect 660 710 760 724
rect 390 646 490 660
rect 390 594 414 646
rect 466 594 490 646
rect 390 580 490 594
rect 130 520 210 530
rect 120 516 220 520
rect 120 464 144 516
rect 196 464 220 516
rect 120 460 220 464
rect 130 450 210 460
<< labels >>
rlabel via1 s 144 464 196 516 4 A
port 1 nsew signal input
rlabel via1 s 414 594 466 646 4 B
port 2 nsew signal input
rlabel via1 s 684 724 736 776 4 Y
port 3 nsew signal output
rlabel metal1 s 110 720 160 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 420 0 540 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 450 720 540 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 820 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 0 820 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 130 450 210 530 1 A
port 1 nsew signal input
rlabel metal2 s 120 460 220 520 1 A
port 1 nsew signal input
rlabel metal1 s 120 460 220 520 1 A
port 1 nsew signal input
rlabel metal2 s 390 580 490 660 1 B
port 2 nsew signal input
rlabel metal1 s 390 590 490 650 1 B
port 2 nsew signal input
rlabel metal2 s 660 710 760 790 1 Y
port 3 nsew signal output
rlabel metal1 s 660 210 710 1060 1 Y
port 3 nsew signal output
rlabel metal1 s 660 710 740 790 1 Y
port 3 nsew signal output
rlabel metal1 s 660 720 760 780 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 820 1270
string GDS_END 36502
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 30992
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
