magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1750858719
transform 1 0 4563 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1750858719
transform 1 0 3891 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1750858719
transform 1 0 400 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1750858719
transform 1 0 1520 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1750858719
transform 1 0 5749 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1750858719
transform 1 0 5973 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1750858719
transform 1 0 1072 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_7
timestamp 1750858719
transform 1 0 848 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_8
timestamp 1750858719
transform 1 0 4787 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_9
timestamp 1750858719
transform 1 0 3667 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_10
timestamp 1750858719
transform 1 0 5525 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_11
timestamp 1750858719
transform 1 0 6197 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_12
timestamp 1750858719
transform 1 0 2929 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_13
timestamp 1750858719
transform 1 0 2257 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_14
timestamp 1750858719
transform 1 0 2705 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_15
timestamp 1750858719
transform 1 0 2481 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_16
timestamp 1750858719
transform 1 0 6421 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_17
timestamp 1750858719
transform 1 0 3153 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_18
timestamp 1750858719
transform 1 0 2033 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_19
timestamp 1750858719
transform 1 0 5301 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_20
timestamp 1750858719
transform 1 0 1296 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_21
timestamp 1750858719
transform 1 0 624 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_22
timestamp 1750858719
transform 1 0 4115 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_23
timestamp 1750858719
transform 1 0 4339 0 1 3151
box 0 0 1 1
use M1_POLY2$$44754988_2_256x8m81  M1_POLY2$$44754988_2_256x8m81_0
timestamp 1750858719
transform 0 -1 7324 -1 0 10090
box 0 0 1 1
use M1_POLY24310590878126_256x8m81  M1_POLY24310590878126_256x8m81_0
timestamp 1750858719
transform 1 0 9070 0 1 9417
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1750858719
transform 1 0 8267 0 1 10062
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1750858719
transform 1 0 8007 0 1 10386
box 0 0 1 1
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_0
timestamp 1750858719
transform -1 0 7291 0 1 10088
box 0 0 1 1
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_1
timestamp 1750858719
transform 1 0 8562 0 1 9367
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1750858719
transform 1 0 8033 0 1 10469
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1750858719
transform 1 0 10229 0 1 9970
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1750858719
transform 1 0 8560 0 1 9721
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1750858719
transform 1 0 9588 0 1 9676
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1750858719
transform 1 0 7374 0 1 9662
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1750858719
transform 1 0 9197 0 1 10519
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1750858719
transform 1 0 7813 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1750858719
transform 1 0 7374 0 1 10576
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_0
timestamp 1750858719
transform -1 0 11659 0 1 3151
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_1
timestamp 1750858719
transform -1 0 11145 0 1 3756
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_2
timestamp 1750858719
transform -1 0 8277 0 1 3555
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_3
timestamp 1750858719
transform -1 0 9968 0 1 3353
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_4
timestamp 1750858719
transform -1 0 9454 0 1 3958
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1750858719
transform 1 0 8211 0 1 10066
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_0
timestamp 1750858719
transform 1 0 8560 0 1 9721
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_1
timestamp 1750858719
transform 1 0 9588 0 1 9676
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_2
timestamp 1750858719
transform 1 0 7374 0 1 9662
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_0
timestamp 1750858719
transform 1 0 9197 0 1 10519
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_1
timestamp 1750858719
transform 1 0 7813 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_2
timestamp 1750858719
transform 1 0 7374 0 1 10576
box 0 0 1 1
use nmos_1p2$$47342636_256x8m81  nmos_1p2$$47342636_256x8m81_0
timestamp 1750858719
transform 1 0 9059 0 1 10236
box -31 0 -30 1
use nmos_5p04310590878160_256x8m81  nmos_5p04310590878160_256x8m81_0
timestamp 1750858719
transform 1 0 7657 0 1 10240
box 0 0 1 1
use nmos_5p04310590878160_256x8m81  nmos_5p04310590878160_256x8m81_1
timestamp 1750858719
transform 1 0 7433 0 1 10240
box 0 0 1 1
use pmos_1p2$$47109164_256x8m81  pmos_1p2$$47109164_256x8m81_0
timestamp 1750858719
transform 1 0 8940 0 1 9519
box -31 0 -30 1
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_0
timestamp 1750858719
transform 1 0 10222 0 1 632
box -20 -633 1762 7970
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_1
timestamp 1750858719
transform 1 0 6841 0 1 632
box -20 -633 1762 7970
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_2
timestamp 1750858719
transform 1 0 8531 0 1 632
box -20 -633 1762 7970
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_0
timestamp 1750858719
transform -1 0 4372 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_1
timestamp 1750858719
transform -1 0 6006 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_2
timestamp 1750858719
transform -1 0 2739 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_3
timestamp 1750858719
transform -1 0 1105 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_4
timestamp 1750858719
transform 1 0 4082 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_5
timestamp 1750858719
transform 1 0 5716 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_6
timestamp 1750858719
transform 1 0 2449 0 1 10644
box 145 -10152 818 -136
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_7
timestamp 1750858719
transform 1 0 815 0 1 10644
box 145 -10152 818 -136
<< properties >>
string GDS_END 1163040
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1153304
<< end >>
