magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 4090 1660
<< nmos >>
rect 190 210 250 380
rect 540 210 600 380
rect 710 210 770 380
rect 820 210 880 380
rect 1170 210 1230 380
rect 1330 210 1390 380
rect 1500 210 1560 380
rect 1610 210 1670 380
rect 1780 210 1840 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2170 210 2230 380
rect 2340 210 2400 380
rect 2690 210 2750 380
rect 3040 210 3100 380
rect 3150 210 3210 380
rect 3320 210 3380 380
rect 3670 210 3730 380
rect 3840 210 3900 380
<< pmos >>
rect 190 1110 250 1450
rect 510 1110 570 1450
rect 680 1110 740 1450
rect 850 1110 910 1450
rect 1170 1110 1230 1450
rect 1330 1110 1390 1450
rect 1500 1110 1560 1450
rect 1610 1110 1670 1450
rect 1780 1110 1840 1450
rect 1890 1110 1950 1450
rect 2060 1110 2120 1450
rect 2170 1110 2230 1450
rect 2340 1110 2400 1450
rect 2690 1110 2750 1450
rect 3010 1110 3070 1450
rect 3180 1110 3240 1450
rect 3350 1110 3410 1450
rect 3670 1110 3730 1450
rect 3840 1110 3900 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 440 318 540 380
rect 440 272 462 318
rect 508 272 540 318
rect 440 210 540 272
rect 600 318 710 380
rect 600 272 632 318
rect 678 272 710 318
rect 600 210 710 272
rect 770 210 820 380
rect 880 318 980 380
rect 880 272 912 318
rect 958 272 980 318
rect 880 210 980 272
rect 1070 318 1170 380
rect 1070 272 1092 318
rect 1138 272 1170 318
rect 1070 210 1170 272
rect 1230 210 1330 380
rect 1390 318 1500 380
rect 1390 272 1422 318
rect 1468 272 1500 318
rect 1390 210 1500 272
rect 1560 210 1610 380
rect 1670 278 1780 380
rect 1670 232 1702 278
rect 1748 232 1780 278
rect 1670 210 1780 232
rect 1840 210 1890 380
rect 1950 318 2060 380
rect 1950 272 1982 318
rect 2028 272 2060 318
rect 1950 210 2060 272
rect 2120 210 2170 380
rect 2230 318 2340 380
rect 2230 272 2262 318
rect 2308 272 2340 318
rect 2230 210 2340 272
rect 2400 318 2500 380
rect 2400 272 2432 318
rect 2478 272 2500 318
rect 2400 210 2500 272
rect 2590 318 2690 380
rect 2590 272 2612 318
rect 2658 272 2690 318
rect 2590 210 2690 272
rect 2750 318 2850 380
rect 2750 272 2782 318
rect 2828 272 2850 318
rect 2750 210 2850 272
rect 2940 318 3040 380
rect 2940 272 2962 318
rect 3008 272 3040 318
rect 2940 210 3040 272
rect 3100 210 3150 380
rect 3210 318 3320 380
rect 3210 272 3242 318
rect 3288 272 3320 318
rect 3210 210 3320 272
rect 3380 318 3480 380
rect 3380 272 3412 318
rect 3458 272 3480 318
rect 3380 210 3480 272
rect 3570 318 3670 380
rect 3570 272 3592 318
rect 3638 272 3670 318
rect 3570 210 3670 272
rect 3730 318 3840 380
rect 3730 272 3762 318
rect 3808 272 3840 318
rect 3730 210 3840 272
rect 3900 318 4000 380
rect 3900 272 3932 318
rect 3978 272 4000 318
rect 3900 210 4000 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 350 1450
rect 250 1163 282 1397
rect 328 1163 350 1397
rect 250 1110 350 1163
rect 410 1397 510 1450
rect 410 1163 432 1397
rect 478 1163 510 1397
rect 410 1110 510 1163
rect 570 1425 680 1450
rect 570 1285 602 1425
rect 648 1285 680 1425
rect 570 1110 680 1285
rect 740 1425 850 1450
rect 740 1285 772 1425
rect 818 1285 850 1425
rect 740 1110 850 1285
rect 910 1425 1010 1450
rect 910 1285 942 1425
rect 988 1285 1010 1425
rect 910 1110 1010 1285
rect 1070 1397 1170 1450
rect 1070 1163 1092 1397
rect 1138 1163 1170 1397
rect 1070 1110 1170 1163
rect 1230 1110 1330 1450
rect 1390 1397 1500 1450
rect 1390 1163 1422 1397
rect 1468 1163 1500 1397
rect 1390 1110 1500 1163
rect 1560 1110 1610 1450
rect 1670 1397 1780 1450
rect 1670 1163 1702 1397
rect 1748 1163 1780 1397
rect 1670 1110 1780 1163
rect 1840 1110 1890 1450
rect 1950 1425 2060 1450
rect 1950 1285 1982 1425
rect 2028 1285 2060 1425
rect 1950 1110 2060 1285
rect 2120 1110 2170 1450
rect 2230 1425 2340 1450
rect 2230 1285 2262 1425
rect 2308 1285 2340 1425
rect 2230 1110 2340 1285
rect 2400 1397 2500 1450
rect 2400 1163 2432 1397
rect 2478 1163 2500 1397
rect 2400 1110 2500 1163
rect 2590 1397 2690 1450
rect 2590 1163 2612 1397
rect 2658 1163 2690 1397
rect 2590 1110 2690 1163
rect 2750 1397 2850 1450
rect 2750 1163 2782 1397
rect 2828 1163 2850 1397
rect 2750 1110 2850 1163
rect 2910 1430 3010 1450
rect 2910 1290 2932 1430
rect 2978 1290 3010 1430
rect 2910 1110 3010 1290
rect 3070 1428 3180 1450
rect 3070 1382 3102 1428
rect 3148 1382 3180 1428
rect 3070 1110 3180 1382
rect 3240 1388 3350 1450
rect 3240 1342 3272 1388
rect 3318 1342 3350 1388
rect 3240 1110 3350 1342
rect 3410 1397 3510 1450
rect 3410 1163 3442 1397
rect 3488 1163 3510 1397
rect 3410 1110 3510 1163
rect 3570 1397 3670 1450
rect 3570 1163 3592 1397
rect 3638 1163 3670 1397
rect 3570 1110 3670 1163
rect 3730 1397 3840 1450
rect 3730 1163 3762 1397
rect 3808 1163 3840 1397
rect 3730 1110 3840 1163
rect 3900 1397 4000 1450
rect 3900 1163 3932 1397
rect 3978 1163 4000 1397
rect 3900 1110 4000 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 462 272 508 318
rect 632 272 678 318
rect 912 272 958 318
rect 1092 272 1138 318
rect 1422 272 1468 318
rect 1702 232 1748 278
rect 1982 272 2028 318
rect 2262 272 2308 318
rect 2432 272 2478 318
rect 2612 272 2658 318
rect 2782 272 2828 318
rect 2962 272 3008 318
rect 3242 272 3288 318
rect 3412 272 3458 318
rect 3592 272 3638 318
rect 3762 272 3808 318
rect 3932 272 3978 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 432 1163 478 1397
rect 602 1285 648 1425
rect 772 1285 818 1425
rect 942 1285 988 1425
rect 1092 1163 1138 1397
rect 1422 1163 1468 1397
rect 1702 1163 1748 1397
rect 1982 1285 2028 1425
rect 2262 1285 2308 1425
rect 2432 1163 2478 1397
rect 2612 1163 2658 1397
rect 2782 1163 2828 1397
rect 2932 1290 2978 1430
rect 3102 1382 3148 1428
rect 3272 1342 3318 1388
rect 3442 1163 3488 1397
rect 3592 1163 3638 1397
rect 3762 1163 3808 1397
rect 3932 1163 3978 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
rect 980 118 1130 140
rect 980 72 1032 118
rect 1078 72 1130 118
rect 980 50 1130 72
rect 1210 118 1360 140
rect 1210 72 1262 118
rect 1308 72 1360 118
rect 1210 50 1360 72
rect 1440 118 1590 140
rect 1440 72 1492 118
rect 1538 72 1590 118
rect 1440 50 1590 72
rect 1670 118 1820 140
rect 1670 72 1722 118
rect 1768 72 1820 118
rect 1670 50 1820 72
rect 1900 118 2050 140
rect 1900 72 1952 118
rect 1998 72 2050 118
rect 1900 50 2050 72
rect 2130 118 2280 140
rect 2130 72 2182 118
rect 2228 72 2280 118
rect 2130 50 2280 72
rect 2360 118 2510 140
rect 2360 72 2412 118
rect 2458 72 2510 118
rect 2360 50 2510 72
rect 2590 118 2740 140
rect 2590 72 2642 118
rect 2688 72 2740 118
rect 2590 50 2740 72
rect 2820 118 2970 140
rect 2820 72 2872 118
rect 2918 72 2970 118
rect 2820 50 2970 72
rect 3050 118 3200 140
rect 3050 72 3102 118
rect 3148 72 3200 118
rect 3050 50 3200 72
rect 3280 118 3430 140
rect 3280 72 3332 118
rect 3378 72 3430 118
rect 3280 50 3430 72
rect 3510 118 3660 140
rect 3510 72 3562 118
rect 3608 72 3660 118
rect 3510 50 3660 72
rect 3740 118 3890 140
rect 3740 72 3792 118
rect 3838 72 3890 118
rect 3740 50 3890 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
rect 980 1588 1130 1610
rect 980 1542 1032 1588
rect 1078 1542 1130 1588
rect 980 1520 1130 1542
rect 1210 1588 1360 1610
rect 1210 1542 1262 1588
rect 1308 1542 1360 1588
rect 1210 1520 1360 1542
rect 1440 1588 1590 1610
rect 1440 1542 1492 1588
rect 1538 1542 1590 1588
rect 1440 1520 1590 1542
rect 1670 1588 1820 1610
rect 1670 1542 1722 1588
rect 1768 1542 1820 1588
rect 1670 1520 1820 1542
rect 1900 1588 2050 1610
rect 1900 1542 1952 1588
rect 1998 1542 2050 1588
rect 1900 1520 2050 1542
rect 2130 1588 2280 1610
rect 2130 1542 2182 1588
rect 2228 1542 2280 1588
rect 2130 1520 2280 1542
rect 2360 1588 2510 1610
rect 2360 1542 2412 1588
rect 2458 1542 2510 1588
rect 2360 1520 2510 1542
rect 2590 1588 2740 1610
rect 2590 1542 2642 1588
rect 2688 1542 2740 1588
rect 2590 1520 2740 1542
rect 2820 1588 2970 1610
rect 2820 1542 2872 1588
rect 2918 1542 2970 1588
rect 2820 1520 2970 1542
rect 3050 1588 3200 1610
rect 3050 1542 3102 1588
rect 3148 1542 3200 1588
rect 3050 1520 3200 1542
rect 3280 1588 3430 1610
rect 3280 1542 3332 1588
rect 3378 1542 3430 1588
rect 3280 1520 3430 1542
rect 3510 1588 3660 1610
rect 3510 1542 3562 1588
rect 3608 1542 3660 1588
rect 3510 1520 3660 1542
rect 3740 1588 3890 1610
rect 3740 1542 3792 1588
rect 3838 1542 3890 1588
rect 3740 1520 3890 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
rect 1032 72 1078 118
rect 1262 72 1308 118
rect 1492 72 1538 118
rect 1722 72 1768 118
rect 1952 72 1998 118
rect 2182 72 2228 118
rect 2412 72 2458 118
rect 2642 72 2688 118
rect 2872 72 2918 118
rect 3102 72 3148 118
rect 3332 72 3378 118
rect 3562 72 3608 118
rect 3792 72 3838 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
rect 1032 1542 1078 1588
rect 1262 1542 1308 1588
rect 1492 1542 1538 1588
rect 1722 1542 1768 1588
rect 1952 1542 1998 1588
rect 2182 1542 2228 1588
rect 2412 1542 2458 1588
rect 2642 1542 2688 1588
rect 2872 1542 2918 1588
rect 3102 1542 3148 1588
rect 3332 1542 3378 1588
rect 3562 1542 3608 1588
rect 3792 1542 3838 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 510 1450 570 1500
rect 680 1450 740 1500
rect 850 1450 910 1500
rect 1170 1450 1230 1500
rect 1330 1450 1390 1500
rect 1500 1450 1560 1500
rect 1610 1450 1670 1500
rect 1780 1450 1840 1500
rect 1890 1450 1950 1500
rect 2060 1450 2120 1500
rect 2170 1450 2230 1500
rect 2340 1450 2400 1500
rect 2690 1450 2750 1500
rect 3010 1450 3070 1500
rect 3180 1450 3240 1500
rect 3350 1450 3410 1500
rect 3670 1450 3730 1500
rect 3840 1450 3900 1500
rect 190 1060 250 1110
rect 120 1038 250 1060
rect 120 992 142 1038
rect 188 992 250 1038
rect 120 970 250 992
rect 190 380 250 970
rect 510 800 570 1110
rect 680 930 740 1110
rect 680 903 800 930
rect 680 857 707 903
rect 753 857 800 903
rect 680 830 800 857
rect 510 773 630 800
rect 510 727 557 773
rect 603 727 630 773
rect 510 700 630 727
rect 510 650 570 700
rect 510 610 600 650
rect 540 380 600 610
rect 680 470 740 830
rect 850 800 910 1110
rect 1170 800 1230 1110
rect 1330 930 1390 1110
rect 1330 903 1430 930
rect 1330 857 1357 903
rect 1403 857 1430 903
rect 1330 830 1430 857
rect 850 773 990 800
rect 850 727 907 773
rect 953 727 990 773
rect 850 700 990 727
rect 1170 773 1290 800
rect 1170 727 1217 773
rect 1263 727 1290 773
rect 1170 700 1290 727
rect 850 470 910 700
rect 680 430 770 470
rect 710 380 770 430
rect 820 430 910 470
rect 820 380 880 430
rect 1170 380 1230 700
rect 1500 660 1560 1110
rect 1610 1060 1670 1110
rect 1780 1060 1840 1110
rect 1610 1033 1840 1060
rect 1610 990 1647 1033
rect 1620 987 1647 990
rect 1693 990 1840 1033
rect 1693 987 1720 990
rect 1620 940 1720 987
rect 1890 660 1950 1110
rect 2060 930 2120 1110
rect 2020 903 2120 930
rect 2020 857 2047 903
rect 2093 857 2120 903
rect 2020 830 2120 857
rect 2170 800 2230 1110
rect 2340 930 2400 1110
rect 2340 903 2440 930
rect 2340 857 2367 903
rect 2413 857 2440 903
rect 2340 830 2440 857
rect 2160 773 2260 800
rect 2160 727 2187 773
rect 2233 727 2260 773
rect 2160 700 2260 727
rect 2020 660 2120 670
rect 1330 643 2120 660
rect 1330 600 2047 643
rect 1330 380 1390 600
rect 2020 597 2047 600
rect 2093 597 2120 643
rect 2020 570 2120 597
rect 1460 513 1560 540
rect 1620 520 1720 540
rect 1460 467 1487 513
rect 1533 467 1560 513
rect 1460 440 1560 467
rect 1500 380 1560 440
rect 1610 513 1840 520
rect 1610 467 1647 513
rect 1693 467 1840 513
rect 1610 440 1840 467
rect 1610 380 1670 440
rect 1780 380 1840 440
rect 1890 503 1990 530
rect 1890 457 1917 503
rect 1963 457 1990 503
rect 1890 430 1990 457
rect 1890 380 1950 430
rect 2060 380 2120 570
rect 2170 380 2230 700
rect 2340 380 2400 830
rect 2690 670 2750 1110
rect 2690 648 2820 670
rect 2690 602 2752 648
rect 2798 602 2820 648
rect 2690 580 2820 602
rect 2690 380 2750 580
rect 3010 530 3070 1110
rect 3180 930 3240 1110
rect 3120 903 3240 930
rect 3120 857 3167 903
rect 3213 857 3240 903
rect 3120 830 3240 857
rect 2930 503 3070 530
rect 2930 457 2967 503
rect 3013 470 3070 503
rect 3180 470 3240 830
rect 3350 650 3410 1110
rect 3670 670 3730 1110
rect 3840 930 3900 1110
rect 3780 903 3900 930
rect 3780 857 3807 903
rect 3853 857 3900 903
rect 3780 830 3900 857
rect 3013 457 3100 470
rect 2930 430 3100 457
rect 3040 380 3100 430
rect 3150 430 3240 470
rect 3320 610 3410 650
rect 3610 643 3730 670
rect 3320 530 3380 610
rect 3610 597 3657 643
rect 3703 597 3730 643
rect 3610 570 3730 597
rect 3320 503 3440 530
rect 3320 457 3367 503
rect 3413 457 3440 503
rect 3320 430 3440 457
rect 3150 380 3210 430
rect 3320 380 3380 430
rect 3670 380 3730 570
rect 3840 380 3900 830
rect 190 160 250 210
rect 540 160 600 210
rect 710 160 770 210
rect 820 160 880 210
rect 1170 160 1230 210
rect 1330 160 1390 210
rect 1500 160 1560 210
rect 1610 160 1670 210
rect 1780 160 1840 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2170 160 2230 210
rect 2340 160 2400 210
rect 2690 160 2750 210
rect 3040 160 3100 210
rect 3150 160 3210 210
rect 3320 160 3380 210
rect 3670 160 3730 210
rect 3840 160 3900 210
<< polycontact >>
rect 142 992 188 1038
rect 707 857 753 903
rect 557 727 603 773
rect 1357 857 1403 903
rect 907 727 953 773
rect 1217 727 1263 773
rect 1647 987 1693 1033
rect 2047 857 2093 903
rect 2367 857 2413 903
rect 2187 727 2233 773
rect 2047 597 2093 643
rect 1487 467 1533 513
rect 1647 467 1693 513
rect 1917 457 1963 503
rect 2752 602 2798 648
rect 3167 857 3213 903
rect 2967 457 3013 503
rect 3807 857 3853 903
rect 3657 597 3703 643
rect 3367 457 3413 503
<< metal1 >>
rect 0 1588 4090 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1032 1588
rect 1078 1542 1262 1588
rect 1308 1542 1492 1588
rect 1538 1542 1722 1588
rect 1768 1542 1952 1588
rect 1998 1542 2182 1588
rect 2228 1542 2412 1588
rect 2458 1542 2642 1588
rect 2688 1542 2872 1588
rect 2918 1542 3102 1588
rect 3148 1542 3332 1588
rect 3378 1542 3562 1588
rect 3608 1542 3792 1588
rect 3838 1542 4090 1588
rect 0 1520 4090 1542
rect 110 1397 160 1520
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1110 160 1163
rect 280 1397 330 1450
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 110 1038 210 1040
rect 110 1036 142 1038
rect 110 984 134 1036
rect 188 992 210 1038
rect 186 984 210 992
rect 110 980 210 984
rect 280 520 330 1163
rect 430 1397 480 1450
rect 430 1163 432 1397
rect 478 1163 480 1397
rect 430 570 480 1163
rect 600 1425 650 1450
rect 600 1285 602 1425
rect 648 1285 650 1425
rect 600 1210 650 1285
rect 770 1425 820 1520
rect 770 1285 772 1425
rect 818 1285 820 1425
rect 770 1260 820 1285
rect 940 1425 990 1450
rect 940 1285 942 1425
rect 988 1285 990 1425
rect 940 1210 990 1285
rect 600 1160 990 1210
rect 1090 1397 1140 1520
rect 1090 1163 1092 1397
rect 1138 1163 1140 1397
rect 1090 1110 1140 1163
rect 1420 1397 1470 1450
rect 1420 1163 1422 1397
rect 1468 1163 1470 1397
rect 1420 1060 1470 1163
rect 1700 1397 1750 1520
rect 1700 1163 1702 1397
rect 1748 1163 1750 1397
rect 1980 1425 2030 1450
rect 1980 1285 1982 1425
rect 2028 1285 2030 1425
rect 1980 1260 2030 1285
rect 2260 1425 2310 1520
rect 2260 1285 2262 1425
rect 2308 1285 2310 1425
rect 2260 1260 2310 1285
rect 2430 1397 2480 1450
rect 1700 1110 1750 1163
rect 1800 1210 2030 1260
rect 1090 1010 1470 1060
rect 1620 1033 1720 1040
rect 680 906 780 910
rect 680 854 704 906
rect 756 854 780 906
rect 680 850 780 854
rect 1090 780 1140 1010
rect 1620 987 1647 1033
rect 1693 987 1720 1033
rect 1620 980 1720 987
rect 1330 906 1560 910
rect 1330 903 1484 906
rect 1330 857 1357 903
rect 1403 857 1484 903
rect 1330 854 1484 857
rect 1536 854 1560 906
rect 1330 850 1560 854
rect 530 776 630 780
rect 530 724 554 776
rect 606 724 630 776
rect 530 720 630 724
rect 880 776 1140 780
rect 880 724 904 776
rect 956 724 1140 776
rect 880 720 1140 724
rect 1190 776 1290 780
rect 1190 724 1214 776
rect 1266 724 1290 776
rect 1190 720 1290 724
rect 430 520 680 570
rect 900 520 950 530
rect 1090 520 1140 720
rect 1480 520 1540 850
rect 1640 520 1700 980
rect 1800 760 1850 1210
rect 2430 1163 2432 1397
rect 2478 1163 2480 1397
rect 2150 1036 2250 1040
rect 2150 984 2174 1036
rect 2226 984 2250 1036
rect 2150 980 2250 984
rect 2430 1020 2480 1163
rect 2610 1397 2660 1450
rect 2610 1163 2612 1397
rect 2658 1163 2660 1397
rect 2610 1130 2660 1163
rect 1790 710 1850 760
rect 1910 906 2120 910
rect 1910 854 2044 906
rect 2096 854 2120 906
rect 1910 850 2120 854
rect 260 516 360 520
rect 260 464 284 516
rect 336 464 360 516
rect 260 460 360 464
rect 630 516 980 520
rect 630 464 904 516
rect 956 464 980 516
rect 1090 470 1290 520
rect 630 460 980 464
rect 280 450 340 460
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 450
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 460 318 510 380
rect 460 272 462 318
rect 508 272 510 318
rect 460 140 510 272
rect 630 318 680 460
rect 900 450 950 460
rect 1210 380 1290 470
rect 1460 513 1560 520
rect 1460 467 1487 513
rect 1533 467 1560 513
rect 1460 460 1560 467
rect 1620 516 1720 520
rect 1620 464 1644 516
rect 1696 464 1720 516
rect 1620 460 1720 464
rect 1790 390 1840 710
rect 1910 510 1970 850
rect 2170 780 2230 980
rect 2430 970 2540 1020
rect 2340 906 2440 910
rect 2340 854 2364 906
rect 2416 854 2440 906
rect 2340 850 2440 854
rect 2490 780 2540 970
rect 2600 910 2660 1130
rect 2780 1397 2830 1520
rect 2780 1163 2782 1397
rect 2828 1163 2830 1397
rect 2930 1430 2980 1450
rect 2930 1290 2932 1430
rect 2978 1310 2980 1430
rect 3100 1428 3150 1520
rect 3100 1382 3102 1428
rect 3148 1382 3150 1428
rect 3100 1360 3150 1382
rect 3270 1388 3320 1450
rect 3270 1342 3272 1388
rect 3318 1342 3320 1388
rect 3270 1310 3320 1342
rect 2978 1290 3320 1310
rect 2930 1260 3320 1290
rect 3440 1397 3490 1450
rect 2780 1110 2830 1163
rect 3440 1163 3442 1397
rect 3488 1163 3490 1397
rect 2960 1040 3020 1060
rect 3440 1040 3490 1163
rect 3590 1397 3640 1450
rect 3590 1163 3592 1397
rect 3638 1163 3640 1397
rect 2960 1036 3520 1040
rect 2960 984 2964 1036
rect 3016 984 3444 1036
rect 3496 984 3520 1036
rect 2960 980 3520 984
rect 2960 960 3020 980
rect 2590 906 2680 910
rect 2590 854 2604 906
rect 2656 854 2680 906
rect 2590 850 2680 854
rect 3140 906 3240 910
rect 3140 854 3164 906
rect 3216 854 3240 906
rect 3140 850 3240 854
rect 2160 776 2260 780
rect 2160 724 2184 776
rect 2236 724 2260 776
rect 2160 720 2260 724
rect 2430 730 2540 780
rect 2020 646 2120 650
rect 2020 594 2044 646
rect 2096 594 2120 646
rect 2020 590 2120 594
rect 2430 646 2490 730
rect 2430 594 2434 646
rect 2486 594 2490 646
rect 2430 570 2490 594
rect 1890 503 1990 510
rect 1890 457 1917 503
rect 1963 457 1990 503
rect 1890 450 1990 457
rect 1790 386 2060 390
rect 630 272 632 318
rect 678 272 680 318
rect 630 210 680 272
rect 910 318 960 380
rect 910 272 912 318
rect 958 272 960 318
rect 910 140 960 272
rect 1090 318 1140 380
rect 1210 330 1470 380
rect 1790 340 1984 386
rect 1090 272 1092 318
rect 1138 272 1140 318
rect 1090 140 1140 272
rect 1420 318 1470 330
rect 1420 272 1422 318
rect 1468 272 1470 318
rect 1980 334 1984 340
rect 2036 334 2060 386
rect 1980 330 2060 334
rect 1980 318 2030 330
rect 1420 210 1470 272
rect 1700 278 1750 300
rect 1700 232 1702 278
rect 1748 232 1750 278
rect 1700 140 1750 232
rect 1980 272 1982 318
rect 2028 272 2030 318
rect 1980 210 2030 272
rect 2260 318 2310 380
rect 2260 272 2262 318
rect 2308 272 2310 318
rect 2260 140 2310 272
rect 2430 318 2480 570
rect 2600 360 2660 850
rect 3440 650 3490 980
rect 3590 910 3640 1163
rect 3760 1397 3810 1520
rect 3760 1163 3762 1397
rect 3808 1163 3810 1397
rect 3760 1110 3810 1163
rect 3930 1397 3980 1450
rect 3930 1163 3932 1397
rect 3978 1163 3980 1397
rect 3930 1050 3980 1163
rect 3930 1036 4030 1050
rect 3930 984 3954 1036
rect 4006 984 4030 1036
rect 3930 980 4030 984
rect 3930 970 4020 980
rect 3590 906 3880 910
rect 3590 854 3804 906
rect 3856 854 3880 906
rect 3590 850 3880 854
rect 2730 648 2830 650
rect 2730 602 2752 648
rect 2798 646 2830 648
rect 2730 594 2754 602
rect 2806 594 2830 646
rect 2730 590 2830 594
rect 3240 646 3730 650
rect 3240 594 3654 646
rect 3706 594 3730 646
rect 3240 590 3730 594
rect 2940 506 3040 510
rect 2940 454 2964 506
rect 3016 454 3040 506
rect 2940 450 3040 454
rect 2430 272 2432 318
rect 2478 272 2480 318
rect 2430 210 2480 272
rect 2610 318 2660 360
rect 2610 272 2612 318
rect 2658 272 2660 318
rect 2610 210 2660 272
rect 2780 318 2830 380
rect 2780 272 2782 318
rect 2828 272 2830 318
rect 2780 140 2830 272
rect 2960 318 3010 380
rect 2960 272 2962 318
rect 3008 272 3010 318
rect 2960 140 3010 272
rect 3240 318 3290 590
rect 3340 506 3440 510
rect 3340 454 3364 506
rect 3416 454 3440 506
rect 3810 480 3860 850
rect 3340 450 3440 454
rect 3590 430 3860 480
rect 3240 272 3242 318
rect 3288 272 3290 318
rect 3240 210 3290 272
rect 3410 318 3460 380
rect 3410 272 3412 318
rect 3458 272 3460 318
rect 3410 140 3460 272
rect 3590 318 3640 430
rect 3590 272 3592 318
rect 3638 272 3640 318
rect 3590 210 3640 272
rect 3760 318 3810 380
rect 3760 272 3762 318
rect 3808 272 3810 318
rect 3760 140 3810 272
rect 3930 318 3980 970
rect 3930 272 3932 318
rect 3978 272 3980 318
rect 3930 210 3980 272
rect 0 118 4090 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1032 118
rect 1078 72 1262 118
rect 1308 72 1492 118
rect 1538 72 1722 118
rect 1768 72 1952 118
rect 1998 72 2182 118
rect 2228 72 2412 118
rect 2458 72 2642 118
rect 2688 72 2872 118
rect 2918 72 3102 118
rect 3148 72 3332 118
rect 3378 72 3562 118
rect 3608 72 3792 118
rect 3838 72 4090 118
rect 0 0 4090 72
<< via1 >>
rect 134 992 142 1036
rect 142 992 186 1036
rect 134 984 186 992
rect 704 903 756 906
rect 704 857 707 903
rect 707 857 753 903
rect 753 857 756 903
rect 704 854 756 857
rect 1484 854 1536 906
rect 554 773 606 776
rect 554 727 557 773
rect 557 727 603 773
rect 603 727 606 773
rect 554 724 606 727
rect 904 773 956 776
rect 904 727 907 773
rect 907 727 953 773
rect 953 727 956 773
rect 904 724 956 727
rect 1214 773 1266 776
rect 1214 727 1217 773
rect 1217 727 1263 773
rect 1263 727 1266 773
rect 1214 724 1266 727
rect 2174 984 2226 1036
rect 2044 903 2096 906
rect 2044 857 2047 903
rect 2047 857 2093 903
rect 2093 857 2096 903
rect 2044 854 2096 857
rect 284 464 336 516
rect 904 464 956 516
rect 1644 513 1696 516
rect 1644 467 1647 513
rect 1647 467 1693 513
rect 1693 467 1696 513
rect 1644 464 1696 467
rect 2364 903 2416 906
rect 2364 857 2367 903
rect 2367 857 2413 903
rect 2413 857 2416 903
rect 2364 854 2416 857
rect 2964 984 3016 1036
rect 3444 984 3496 1036
rect 2604 854 2656 906
rect 3164 903 3216 906
rect 3164 857 3167 903
rect 3167 857 3213 903
rect 3213 857 3216 903
rect 3164 854 3216 857
rect 2184 773 2236 776
rect 2184 727 2187 773
rect 2187 727 2233 773
rect 2233 727 2236 773
rect 2184 724 2236 727
rect 2044 643 2096 646
rect 2044 597 2047 643
rect 2047 597 2093 643
rect 2093 597 2096 643
rect 2044 594 2096 597
rect 2434 594 2486 646
rect 1984 334 2036 386
rect 3954 984 4006 1036
rect 3804 903 3856 906
rect 3804 857 3807 903
rect 3807 857 3853 903
rect 3853 857 3856 903
rect 3804 854 3856 857
rect 2754 602 2798 646
rect 2798 602 2806 646
rect 2754 594 2806 602
rect 3654 643 3706 646
rect 3654 597 3657 643
rect 3657 597 3703 643
rect 3703 597 3706 643
rect 3654 594 3706 597
rect 2964 503 3016 506
rect 2964 457 2967 503
rect 2967 457 3013 503
rect 3013 457 3016 503
rect 2964 454 3016 457
rect 3364 503 3416 506
rect 3364 457 3367 503
rect 3367 457 3413 503
rect 3413 457 3416 503
rect 3364 454 3416 457
<< metal2 >>
rect 700 1110 3220 1170
rect 110 1036 210 1050
rect 110 984 134 1036
rect 186 984 210 1036
rect 110 970 210 984
rect 700 920 760 1110
rect 2160 1040 2240 1050
rect 2950 1040 3030 1050
rect 2150 1036 3040 1040
rect 2150 984 2174 1036
rect 2226 984 2964 1036
rect 3016 984 3040 1036
rect 2150 980 3040 984
rect 2160 970 2240 980
rect 2950 970 3030 980
rect 3160 920 3220 1110
rect 3420 1036 3520 1050
rect 3940 1040 4020 1050
rect 3420 984 3444 1036
rect 3496 984 3520 1036
rect 3420 970 3520 984
rect 3930 1036 4030 1040
rect 3930 984 3954 1036
rect 4006 984 4030 1036
rect 3930 980 4030 984
rect 3940 970 4020 980
rect 680 906 780 920
rect 680 854 704 906
rect 756 854 780 906
rect 680 840 780 854
rect 1460 910 1550 920
rect 2020 910 2120 920
rect 2350 910 2430 920
rect 2590 910 2680 920
rect 1460 906 2680 910
rect 1460 854 1484 906
rect 1536 854 2044 906
rect 2096 854 2364 906
rect 2416 854 2604 906
rect 2656 854 2680 906
rect 1460 850 2680 854
rect 1460 840 1550 850
rect 2020 840 2120 850
rect 2350 840 2430 850
rect 2590 840 2680 850
rect 3140 906 3240 920
rect 3790 910 3870 920
rect 3140 854 3164 906
rect 3216 854 3240 906
rect 3140 840 3240 854
rect 3780 906 3880 910
rect 3780 854 3804 906
rect 3856 854 3880 906
rect 3780 850 3880 854
rect 3790 840 3870 850
rect 530 776 630 790
rect 530 724 554 776
rect 606 724 630 776
rect 530 710 630 724
rect 880 776 980 790
rect 880 724 904 776
rect 956 724 980 776
rect 880 710 980 724
rect 1190 776 1290 790
rect 2170 780 2250 790
rect 1190 724 1214 776
rect 1266 724 1290 776
rect 1190 710 1290 724
rect 2160 776 2260 780
rect 2160 724 2184 776
rect 2236 724 2260 776
rect 2160 720 2260 724
rect 2170 710 2250 720
rect 260 520 360 530
rect 550 520 610 710
rect 2030 650 2110 660
rect 2420 650 2500 660
rect 2020 646 2520 650
rect 2020 594 2044 646
rect 2096 594 2434 646
rect 2486 594 2520 646
rect 2020 590 2520 594
rect 2730 646 2830 660
rect 3640 650 3720 660
rect 2730 594 2754 646
rect 2806 594 2830 646
rect 2030 580 2110 590
rect 2420 580 2500 590
rect 2730 580 2830 594
rect 3570 646 3730 650
rect 3570 594 3654 646
rect 3706 594 3730 646
rect 3570 590 3730 594
rect 3640 580 3720 590
rect 260 516 610 520
rect 260 464 284 516
rect 336 464 610 516
rect 260 460 610 464
rect 260 450 360 460
rect 550 260 610 460
rect 880 520 980 530
rect 1630 520 1710 530
rect 880 516 1720 520
rect 880 464 904 516
rect 956 464 1644 516
rect 1696 464 1720 516
rect 880 460 1720 464
rect 2940 506 3040 520
rect 880 450 980 460
rect 1630 450 1710 460
rect 2940 454 2964 506
rect 3016 454 3040 506
rect 2940 440 3040 454
rect 3320 506 3440 520
rect 3320 454 3364 506
rect 3416 454 3440 506
rect 3320 440 3440 454
rect 1970 390 2050 400
rect 2940 390 3020 440
rect 1960 386 3020 390
rect 1960 334 1984 386
rect 2036 334 3020 386
rect 1960 330 3020 334
rect 1970 320 2050 330
rect 3320 260 3380 440
rect 550 200 3380 260
<< labels >>
rlabel via1 s 1214 724 1266 776 4 D
port 1 nsew signal input
rlabel via1 s 3954 984 4006 1036 4 Q
port 2 nsew signal output
rlabel via1 s 3804 854 3856 906 4 QN
port 3 nsew signal output
rlabel via1 s 2754 594 2806 646 4 CLK
port 4 nsew clock input
rlabel via1 s 134 984 186 1036 4 RN
port 5 nsew signal input
rlabel via1 s 3164 854 3216 906 4 SN
port 6 nsew signal output
rlabel metal1 s 110 1110 160 1660 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 770 1260 820 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1090 1110 1140 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1700 1110 1750 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2260 1260 2310 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2780 1110 2830 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3100 1360 3150 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3760 1110 3810 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 1520 4090 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 460 0 510 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 910 0 960 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1090 0 1140 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1700 0 1750 300 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2260 0 2310 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2780 0 2830 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2960 0 3010 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3410 0 3460 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3760 0 3810 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 0 4090 140 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal2 s 2730 580 2830 660 1 CLK
port 4 nsew clock input
rlabel metal1 s 2730 590 2830 650 1 CLK
port 4 nsew clock input
rlabel metal2 s 1190 710 1290 790 1 D
port 1 nsew signal input
rlabel metal1 s 1190 720 1290 780 1 D
port 1 nsew signal input
rlabel metal2 s 3940 970 4020 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3930 980 4030 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 3930 210 3980 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 3930 970 4020 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 3930 980 4030 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3790 840 3870 920 1 QN
port 3 nsew signal output
rlabel metal2 s 3780 850 3880 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 210 3640 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 850 3640 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 430 3860 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3810 430 3860 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 850 3880 910 1 QN
port 3 nsew signal output
rlabel metal2 s 110 970 210 1050 1 RN
port 5 nsew signal input
rlabel metal1 s 110 980 210 1040 1 RN
port 5 nsew signal input
rlabel via1 s 704 854 756 906 1 SN
port 6 nsew signal output
rlabel metal2 s 700 840 760 1170 1 SN
port 6 nsew signal output
rlabel metal2 s 680 840 780 920 1 SN
port 6 nsew signal output
rlabel metal2 s 3160 840 3220 1170 1 SN
port 6 nsew signal output
rlabel metal2 s 700 1110 3220 1170 1 SN
port 6 nsew signal output
rlabel metal2 s 3140 840 3240 920 1 SN
port 6 nsew signal output
rlabel metal1 s 680 850 780 910 1 SN
port 6 nsew signal output
rlabel metal1 s 3140 850 3240 910 1 SN
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 4090 1660
string GDS_END 375160
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 344958
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
