magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< obsm1 >>
rect -32 13108 15032 69957
<< metal2 >>
rect 272 69069 2172 70000
rect 2752 69069 4802 70000
rect 5122 69069 7172 70000
rect 7828 69069 9878 70000
rect 10198 69069 12248 70000
rect 12828 69069 14728 70000
<< obsm2 >>
rect 0 69009 212 69678
rect 2232 69009 2692 69678
rect 4862 69009 5062 69678
rect 7232 69009 7768 69678
rect 9938 69009 10138 69678
rect 12308 69009 12768 69678
rect 14788 69009 15000 69678
rect 0 0 15000 69009
<< metal3 >>
rect 0 68400 2502 69678
rect 0 66800 326 68200
rect 12498 68400 15000 69678
rect 0 65200 2502 66600
rect 0 63600 200 65000
rect 14674 66800 15000 68200
rect 12498 65200 15000 66600
rect 0 62000 326 63400
rect 14800 63600 15000 65000
rect 0 60400 2502 61800
rect 0 58800 326 60200
rect 14674 62000 15000 63400
rect 12498 60400 15000 61800
rect 0 57200 2502 58600
rect 0 55600 326 57000
rect 14674 58800 15000 60200
rect 12498 57200 15000 58600
rect 0 54000 326 55400
rect 0 52400 326 53800
rect 0 50800 326 52200
rect 0 49200 200 50600
rect 14674 55600 15000 57000
rect 14674 54000 15000 55400
rect 14674 52400 15000 53800
rect 14674 50800 15000 52200
rect 0 46000 2502 49000
rect 0 42800 326 45800
rect 14800 49200 15000 50600
rect 12498 46000 15000 49000
rect 0 41200 326 42600
rect 14674 42800 15000 45800
rect 0 39600 2502 41000
rect 0 36400 326 39400
rect 14674 41200 15000 42600
rect 12498 39600 15000 41000
rect 0 33200 326 36200
rect 0 30000 326 33000
rect 0 26800 326 29800
rect 14674 36400 15000 39400
rect 14674 33200 15000 36200
rect 14674 30000 15000 33000
rect 0 25200 2502 26600
rect 0 23600 326 25000
rect 14674 26800 15000 29800
rect 12498 25200 15000 26600
rect 0 20400 2502 23400
rect 0 17200 2502 20200
rect 0 14000 2502 17000
rect 14674 23600 15000 25000
rect 12498 20400 15000 23400
rect 12498 17200 15000 20200
rect 12498 14000 15000 17000
<< obsm3 >>
rect 2862 68040 12138 69678
rect 686 66960 14314 68040
rect 2862 64840 12138 66960
rect 560 63760 14440 64840
rect 686 62160 14314 63760
rect 2862 60040 12138 62160
rect 686 58960 14314 60040
rect 2862 56840 12138 58960
rect 686 50440 14314 56840
rect 560 49360 14440 50440
rect 2862 45640 12138 49360
rect 686 41360 14314 45640
rect 2862 39240 12138 41360
rect 686 26960 14314 39240
rect 2862 24840 12138 26960
rect 686 23760 14314 24840
rect 2862 13640 12138 23760
rect 200 0 14800 13640
<< labels >>
rlabel metal3 s 14674 23600 15000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 36400 15000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 33200 15000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 30000 15000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 26800 15000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 42800 15000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 41200 15000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 50800 15000 52200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 55600 15000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 54000 15000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 52400 15000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 58800 15000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 62000 15000 63400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14674 66800 15000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 272 69069 2172 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 2752 69069 4802 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 5122 69069 7172 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 7828 69069 9878 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 10198 69069 12248 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 66800 326 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 62000 326 63400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 326 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 326 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 326 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 326 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 50800 326 52200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 326 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 326 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 326 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 326 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 326 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 326 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 326 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal2 s 12828 69069 14728 70000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 20400 15000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 17200 15000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 14000 15000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 25200 15000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 39600 15000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 46000 15000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 57200 15000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 60400 15000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 65200 15000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 12498 68400 15000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 68400 2502 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 2502 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 2502 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 2502 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 2502 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 2502 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 2502 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 2502 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 2502 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 2502 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 49200 15000 50600 6 VSS
port 3 nsew ground bidirectional
rlabel metal3 s 14800 63600 15000 65000 6 VSS
port 3 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 6 VSS
port 3 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 6 VSS
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD POWER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4039472
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4037764
<< end >>
