magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 960 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
rect 700 720 760 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 318 530 380
rect 420 272 452 318
rect 498 272 530 318
rect 420 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 318 860 380
rect 760 272 792 318
rect 838 272 860 318
rect 760 210 860 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 360 1060
rect 250 773 282 1007
rect 328 773 360 1007
rect 250 720 360 773
rect 420 1007 530 1060
rect 420 773 452 1007
rect 498 773 530 1007
rect 420 720 530 773
rect 590 1007 700 1060
rect 590 773 622 1007
rect 668 773 700 1007
rect 590 720 700 773
rect 760 1007 870 1060
rect 760 773 802 1007
rect 848 773 870 1007
rect 760 720 870 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 792 272 838 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 452 773 498 1007
rect 622 773 668 1007
rect 802 773 848 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 700 1060 760 1110
rect 190 670 250 720
rect 360 670 420 720
rect 530 670 590 720
rect 700 670 760 720
rect 190 620 760 670
rect 190 540 250 620
rect 90 518 250 540
rect 90 472 112 518
rect 158 480 250 518
rect 158 472 760 480
rect 90 450 760 472
rect 190 420 760 450
rect 190 380 250 420
rect 360 380 420 420
rect 530 380 590 420
rect 700 380 760 420
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
<< polycontact >>
rect 112 472 158 518
<< metal1 >>
rect 0 1198 960 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 960 1198
rect 0 1130 960 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 670 330 773
rect 450 1007 500 1130
rect 450 773 452 1007
rect 498 773 500 1007
rect 450 720 500 773
rect 620 1007 670 1060
rect 620 773 622 1007
rect 668 780 670 1007
rect 800 1007 850 1130
rect 668 776 750 780
rect 668 773 674 776
rect 620 724 674 773
rect 726 724 750 776
rect 620 720 750 724
rect 800 773 802 1007
rect 848 773 850 1007
rect 800 720 850 773
rect 620 670 670 720
rect 280 620 670 670
rect 80 518 180 520
rect 80 516 112 518
rect 80 464 104 516
rect 158 472 180 518
rect 156 464 180 472
rect 80 460 180 464
rect 280 480 330 620
rect 620 480 670 620
rect 280 430 670 480
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 430
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 450 318 500 380
rect 450 272 452 318
rect 498 272 500 318
rect 450 140 500 272
rect 620 318 670 430
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 790 318 840 380
rect 790 272 792 318
rect 838 272 840 318
rect 790 140 840 272
rect 0 118 960 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 960 118
rect 0 0 960 72
<< via1 >>
rect 674 724 726 776
rect 104 472 112 516
rect 112 472 156 516
rect 104 464 156 472
<< metal2 >>
rect 660 780 740 790
rect 650 776 750 780
rect 650 724 674 776
rect 726 724 750 776
rect 650 720 750 724
rect 660 710 740 720
rect 80 516 180 530
rect 80 464 104 516
rect 156 464 180 516
rect 80 450 180 464
<< labels >>
rlabel via1 s 104 464 156 516 4 A
port 1 nsew signal input
rlabel via1 s 674 724 726 776 4 Y
port 2 nsew signal output
rlabel metal1 s 110 720 160 1270 4 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 450 720 500 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 800 720 850 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 1130 960 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 450 0 500 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 790 0 840 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 0 960 140 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal2 s 80 450 180 530 1 A
port 1 nsew signal input
rlabel metal1 s 80 460 180 520 1 A
port 1 nsew signal input
rlabel metal2 s 660 710 740 790 1 Y
port 2 nsew signal output
rlabel metal2 s 650 720 750 780 1 Y
port 2 nsew signal output
rlabel metal1 s 280 210 330 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 280 430 670 480 1 Y
port 2 nsew signal output
rlabel metal1 s 280 620 670 670 1 Y
port 2 nsew signal output
rlabel metal1 s 620 210 670 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 620 720 750 780 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 960 1270
string GDS_END 151340
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 145676
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
