magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 5350 870
<< pwell >>
rect -86 -86 5350 352
<< mvnmos >>
rect 124 68 244 232
rect 308 68 428 232
rect 532 68 652 232
rect 716 68 836 232
rect 940 68 1060 232
rect 1124 68 1244 232
rect 1348 68 1468 232
rect 1532 68 1652 232
rect 1890 68 2010 232
rect 2084 68 2204 232
rect 2308 68 2428 232
rect 2492 68 2612 232
rect 2716 68 2836 232
rect 2900 68 3020 232
rect 3124 68 3244 232
rect 3308 68 3428 232
rect 3532 68 3652 232
rect 3716 68 3836 232
rect 3940 68 4060 232
rect 4124 68 4244 232
rect 4348 68 4468 232
rect 4532 68 4652 232
rect 4756 68 4876 232
rect 4940 68 5060 232
<< mvpmos >>
rect 124 472 224 716
rect 328 472 428 716
rect 532 472 632 716
rect 736 472 836 716
rect 940 472 1040 716
rect 1144 472 1244 716
rect 1348 472 1448 716
rect 1552 472 1652 716
rect 1900 472 2000 716
rect 2104 472 2204 716
rect 2308 472 2408 716
rect 2512 472 2612 716
rect 2716 472 2816 716
rect 2920 472 3020 716
rect 3124 472 3224 716
rect 3328 472 3428 716
rect 3532 472 3632 716
rect 3736 472 3836 716
rect 3940 472 4040 716
rect 4144 472 4244 716
rect 4348 472 4448 716
rect 4552 472 4652 716
rect 4756 472 4856 716
rect 4960 472 5060 716
<< mvndiff >>
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 68 308 232
rect 428 127 532 232
rect 428 81 457 127
rect 503 81 532 127
rect 428 68 532 81
rect 652 68 716 232
rect 836 219 940 232
rect 836 173 865 219
rect 911 173 940 219
rect 836 68 940 173
rect 1060 68 1124 232
rect 1244 127 1348 232
rect 1244 81 1273 127
rect 1319 81 1348 127
rect 1244 68 1348 81
rect 1468 68 1532 232
rect 1652 219 1890 232
rect 1652 173 1681 219
rect 1727 173 1815 219
rect 1861 173 1890 219
rect 1652 68 1890 173
rect 2010 68 2084 232
rect 2204 127 2308 232
rect 2204 81 2233 127
rect 2279 81 2308 127
rect 2204 68 2308 81
rect 2428 68 2492 232
rect 2612 219 2716 232
rect 2612 173 2641 219
rect 2687 173 2716 219
rect 2612 68 2716 173
rect 2836 68 2900 232
rect 3020 127 3124 232
rect 3020 81 3049 127
rect 3095 81 3124 127
rect 3020 68 3124 81
rect 3244 68 3308 232
rect 3428 160 3532 232
rect 3428 114 3457 160
rect 3503 114 3532 160
rect 3428 68 3532 114
rect 3652 68 3716 232
rect 3836 127 3940 232
rect 3836 81 3865 127
rect 3911 81 3940 127
rect 3836 68 3940 81
rect 4060 68 4124 232
rect 4244 152 4348 232
rect 4244 106 4273 152
rect 4319 106 4348 152
rect 4244 68 4348 106
rect 4468 68 4532 232
rect 4652 127 4756 232
rect 4652 81 4681 127
rect 4727 81 4756 127
rect 4652 68 4756 81
rect 4876 68 4940 232
rect 5060 219 5148 232
rect 5060 173 5089 219
rect 5135 173 5148 219
rect 5060 68 5148 173
<< mvpdiff >>
rect 36 665 124 716
rect 36 525 49 665
rect 95 525 124 665
rect 36 472 124 525
rect 224 665 328 716
rect 224 525 253 665
rect 299 525 328 665
rect 224 472 328 525
rect 428 665 532 716
rect 428 619 457 665
rect 503 619 532 665
rect 428 472 532 619
rect 632 665 736 716
rect 632 525 661 665
rect 707 525 736 665
rect 632 472 736 525
rect 836 665 940 716
rect 836 619 865 665
rect 911 619 940 665
rect 836 472 940 619
rect 1040 665 1144 716
rect 1040 525 1069 665
rect 1115 525 1144 665
rect 1040 472 1144 525
rect 1244 665 1348 716
rect 1244 619 1273 665
rect 1319 619 1348 665
rect 1244 472 1348 619
rect 1448 665 1552 716
rect 1448 525 1477 665
rect 1523 525 1552 665
rect 1448 472 1552 525
rect 1652 665 1740 716
rect 1652 619 1681 665
rect 1727 619 1740 665
rect 1652 472 1740 619
rect 1812 678 1900 716
rect 1812 632 1825 678
rect 1871 632 1900 678
rect 1812 472 1900 632
rect 2000 552 2104 716
rect 2000 506 2029 552
rect 2075 506 2104 552
rect 2000 472 2104 506
rect 2204 678 2308 716
rect 2204 632 2233 678
rect 2279 632 2308 678
rect 2204 472 2308 632
rect 2408 552 2512 716
rect 2408 506 2437 552
rect 2483 506 2512 552
rect 2408 472 2512 506
rect 2612 678 2716 716
rect 2612 632 2641 678
rect 2687 632 2716 678
rect 2612 472 2716 632
rect 2816 552 2920 716
rect 2816 506 2845 552
rect 2891 506 2920 552
rect 2816 472 2920 506
rect 3020 678 3124 716
rect 3020 632 3049 678
rect 3095 632 3124 678
rect 3020 472 3124 632
rect 3224 552 3328 716
rect 3224 506 3253 552
rect 3299 506 3328 552
rect 3224 472 3328 506
rect 3428 678 3532 716
rect 3428 632 3457 678
rect 3503 632 3532 678
rect 3428 472 3532 632
rect 3632 567 3736 716
rect 3632 521 3661 567
rect 3707 521 3736 567
rect 3632 472 3736 521
rect 3836 678 3940 716
rect 3836 632 3865 678
rect 3911 632 3940 678
rect 3836 472 3940 632
rect 4040 567 4144 716
rect 4040 521 4069 567
rect 4115 521 4144 567
rect 4040 472 4144 521
rect 4244 678 4348 716
rect 4244 632 4273 678
rect 4319 632 4348 678
rect 4244 472 4348 632
rect 4448 567 4552 716
rect 4448 521 4477 567
rect 4523 521 4552 567
rect 4448 472 4552 521
rect 4652 678 4756 716
rect 4652 632 4681 678
rect 4727 632 4756 678
rect 4652 472 4756 632
rect 4856 567 4960 716
rect 4856 521 4885 567
rect 4931 521 4960 567
rect 4856 472 4960 521
rect 5060 665 5148 716
rect 5060 525 5089 665
rect 5135 525 5148 665
rect 5060 472 5148 525
<< mvndiffc >>
rect 49 173 95 219
rect 457 81 503 127
rect 865 173 911 219
rect 1273 81 1319 127
rect 1681 173 1727 219
rect 1815 173 1861 219
rect 2233 81 2279 127
rect 2641 173 2687 219
rect 3049 81 3095 127
rect 3457 114 3503 160
rect 3865 81 3911 127
rect 4273 106 4319 152
rect 4681 81 4727 127
rect 5089 173 5135 219
<< mvpdiffc >>
rect 49 525 95 665
rect 253 525 299 665
rect 457 619 503 665
rect 661 525 707 665
rect 865 619 911 665
rect 1069 525 1115 665
rect 1273 619 1319 665
rect 1477 525 1523 665
rect 1681 619 1727 665
rect 1825 632 1871 678
rect 2029 506 2075 552
rect 2233 632 2279 678
rect 2437 506 2483 552
rect 2641 632 2687 678
rect 2845 506 2891 552
rect 3049 632 3095 678
rect 3253 506 3299 552
rect 3457 632 3503 678
rect 3661 521 3707 567
rect 3865 632 3911 678
rect 4069 521 4115 567
rect 4273 632 4319 678
rect 4477 521 4523 567
rect 4681 632 4727 678
rect 4885 521 4931 567
rect 5089 525 5135 665
<< polysilicon >>
rect 124 716 224 760
rect 328 716 428 760
rect 532 716 632 760
rect 736 716 836 760
rect 940 716 1040 760
rect 1144 716 1244 760
rect 1348 716 1448 760
rect 1552 716 1652 760
rect 1900 716 2000 760
rect 2104 716 2204 760
rect 2308 716 2408 760
rect 2512 716 2612 760
rect 2716 716 2816 760
rect 2920 716 3020 760
rect 3124 716 3224 760
rect 3328 716 3428 760
rect 3532 716 3632 760
rect 3736 716 3836 760
rect 3940 716 4040 760
rect 4144 716 4244 760
rect 4348 716 4448 760
rect 4552 716 4652 760
rect 4756 716 4856 760
rect 4960 716 5060 760
rect 124 313 224 472
rect 124 267 165 313
rect 211 288 224 313
rect 328 415 428 472
rect 328 369 353 415
rect 399 394 428 415
rect 532 415 632 472
rect 532 394 560 415
rect 399 369 560 394
rect 606 369 632 415
rect 328 348 632 369
rect 328 288 428 348
rect 211 267 244 288
rect 124 232 244 267
rect 308 232 428 288
rect 532 288 632 348
rect 736 394 836 472
rect 940 394 1040 472
rect 736 348 1040 394
rect 736 313 836 348
rect 736 288 761 313
rect 532 232 652 288
rect 716 267 761 288
rect 807 267 836 313
rect 716 232 836 267
rect 940 288 1040 348
rect 1144 415 1244 472
rect 1144 369 1169 415
rect 1215 394 1244 415
rect 1348 415 1448 472
rect 1348 394 1361 415
rect 1215 369 1361 394
rect 1407 369 1448 415
rect 1144 348 1448 369
rect 1144 288 1244 348
rect 940 232 1060 288
rect 1124 232 1244 288
rect 1348 288 1448 348
rect 1552 415 1652 472
rect 1552 369 1565 415
rect 1611 369 1652 415
rect 1552 288 1652 369
rect 1900 415 2000 472
rect 1900 369 1937 415
rect 1983 369 2000 415
rect 1900 288 2000 369
rect 2104 414 2204 472
rect 2104 368 2133 414
rect 2179 394 2204 414
rect 2308 414 2408 472
rect 2308 394 2340 414
rect 2179 368 2340 394
rect 2386 368 2408 414
rect 2104 348 2408 368
rect 2104 288 2204 348
rect 1348 232 1468 288
rect 1532 232 1652 288
rect 1890 232 2010 288
rect 2084 232 2204 288
rect 2308 288 2408 348
rect 2512 394 2612 472
rect 2716 394 2816 472
rect 2512 348 2816 394
rect 2512 313 2612 348
rect 2512 288 2535 313
rect 2308 232 2428 288
rect 2492 267 2535 288
rect 2581 267 2612 313
rect 2492 232 2612 267
rect 2716 313 2816 348
rect 2716 267 2745 313
rect 2791 288 2816 313
rect 2920 415 3020 472
rect 2920 369 2945 415
rect 2991 394 3020 415
rect 3124 415 3224 472
rect 3124 394 3148 415
rect 2991 369 3148 394
rect 3194 369 3224 415
rect 3328 407 3428 472
rect 2920 348 3224 369
rect 2920 288 3020 348
rect 2791 267 2836 288
rect 2716 232 2836 267
rect 2900 232 3020 288
rect 3124 288 3224 348
rect 3308 394 3428 407
rect 3308 348 3321 394
rect 3367 348 3428 394
rect 3124 232 3244 288
rect 3308 232 3428 348
rect 3532 439 3632 472
rect 3532 393 3573 439
rect 3619 393 3632 439
rect 3532 288 3632 393
rect 3736 394 3836 472
rect 3940 394 4040 472
rect 3736 348 4040 394
rect 3736 317 3836 348
rect 3736 288 3758 317
rect 3532 232 3652 288
rect 3716 271 3758 288
rect 3804 271 3836 317
rect 3716 232 3836 271
rect 3940 317 4040 348
rect 3940 271 3973 317
rect 4019 288 4040 317
rect 4144 439 4244 472
rect 4144 393 4168 439
rect 4214 394 4244 439
rect 4348 439 4448 472
rect 4348 394 4373 439
rect 4214 393 4373 394
rect 4419 393 4448 439
rect 4144 348 4448 393
rect 4144 288 4244 348
rect 4019 271 4060 288
rect 3940 232 4060 271
rect 4124 232 4244 288
rect 4348 288 4448 348
rect 4552 394 4652 472
rect 4756 394 4856 472
rect 4552 348 4856 394
rect 4552 311 4652 348
rect 4552 288 4565 311
rect 4348 232 4468 288
rect 4532 265 4565 288
rect 4611 265 4652 311
rect 4532 232 4652 265
rect 4756 288 4856 348
rect 4960 439 5060 472
rect 4960 393 4973 439
rect 5019 393 5060 439
rect 4960 288 5060 393
rect 4756 232 4876 288
rect 4940 232 5060 288
rect 124 24 244 68
rect 308 24 428 68
rect 532 24 652 68
rect 716 24 836 68
rect 940 24 1060 68
rect 1124 24 1244 68
rect 1348 24 1468 68
rect 1532 24 1652 68
rect 1890 24 2010 68
rect 2084 24 2204 68
rect 2308 24 2428 68
rect 2492 24 2612 68
rect 2716 24 2836 68
rect 2900 24 3020 68
rect 3124 24 3244 68
rect 3308 24 3428 68
rect 3532 24 3652 68
rect 3716 24 3836 68
rect 3940 24 4060 68
rect 4124 24 4244 68
rect 4348 24 4468 68
rect 4532 24 4652 68
rect 4756 24 4876 68
rect 4940 24 5060 68
<< polycontact >>
rect 165 267 211 313
rect 353 369 399 415
rect 560 369 606 415
rect 761 267 807 313
rect 1169 369 1215 415
rect 1361 369 1407 415
rect 1565 369 1611 415
rect 1937 369 1983 415
rect 2133 368 2179 414
rect 2340 368 2386 414
rect 2535 267 2581 313
rect 2745 267 2791 313
rect 2945 369 2991 415
rect 3148 369 3194 415
rect 3321 348 3367 394
rect 3573 393 3619 439
rect 3758 271 3804 317
rect 3973 271 4019 317
rect 4168 393 4214 439
rect 4373 393 4419 439
rect 4565 265 4611 311
rect 4973 393 5019 439
<< metal1 >>
rect 0 724 5264 844
rect 38 665 106 724
rect 38 525 49 665
rect 95 525 106 665
rect 38 511 106 525
rect 242 665 310 676
rect 242 525 253 665
rect 299 552 310 665
rect 446 665 515 724
rect 446 619 457 665
rect 503 619 515 665
rect 446 608 515 619
rect 650 665 718 676
rect 650 552 661 665
rect 299 525 661 552
rect 707 552 718 665
rect 854 665 922 724
rect 854 619 865 665
rect 911 619 922 665
rect 854 608 922 619
rect 1058 665 1126 676
rect 1058 552 1069 665
rect 707 525 1069 552
rect 1115 552 1126 665
rect 1262 665 1330 724
rect 1262 619 1273 665
rect 1319 619 1330 665
rect 1262 608 1330 619
rect 1466 665 1534 676
rect 1466 552 1477 665
rect 1115 525 1477 552
rect 1523 552 1534 665
rect 1670 665 1738 724
rect 1670 619 1681 665
rect 1727 619 1738 665
rect 1814 632 1825 678
rect 1871 632 2233 678
rect 2279 632 2641 678
rect 2687 632 3049 678
rect 3095 632 3457 678
rect 3503 632 3865 678
rect 3911 632 4273 678
rect 4319 632 4681 678
rect 4727 665 5146 678
rect 4727 632 5089 665
rect 1670 608 1738 619
rect 1523 525 2029 552
rect 242 506 2029 525
rect 2075 506 2437 552
rect 2483 506 2845 552
rect 2891 506 3253 552
rect 3299 506 3310 552
rect 3415 521 3661 567
rect 3707 521 4069 567
rect 4115 521 4477 567
rect 4523 521 4885 567
rect 4931 521 4942 567
rect 5078 525 5089 632
rect 5135 525 5146 665
rect 117 415 1418 424
rect 117 369 353 415
rect 399 369 560 415
rect 606 369 1169 415
rect 1215 369 1361 415
rect 1407 369 1418 415
rect 117 360 1418 369
rect 1464 415 1703 430
rect 1464 369 1565 415
rect 1611 369 1703 415
rect 1464 352 1703 369
rect 1789 415 2032 430
rect 1789 369 1937 415
rect 1983 369 2032 415
rect 1464 313 1524 352
rect 142 267 165 313
rect 211 267 761 313
rect 807 267 1524 313
rect 1789 313 2032 369
rect 2083 415 3251 424
rect 2083 414 2945 415
rect 2083 368 2133 414
rect 2179 368 2340 414
rect 2386 369 2945 414
rect 2991 369 3148 415
rect 3194 369 3251 415
rect 2386 368 3251 369
rect 2083 360 3251 368
rect 3321 394 3367 405
rect 3321 313 3367 348
rect 1789 267 2535 313
rect 2581 267 2745 313
rect 2791 267 3367 313
rect 1126 219 1407 220
rect 38 173 49 219
rect 95 173 865 219
rect 911 174 1681 219
rect 911 173 1172 174
rect 1361 173 1681 174
rect 1727 173 1815 219
rect 1861 173 2641 219
rect 2687 173 3208 219
rect 3162 160 3208 173
rect 3415 160 3461 521
rect 5078 511 5146 525
rect 3556 393 3573 439
rect 3619 393 4168 439
rect 4214 393 4373 439
rect 4419 393 4973 439
rect 5019 393 5134 439
rect 4722 354 5134 393
rect 3507 317 4622 323
rect 3507 271 3758 317
rect 3804 271 3973 317
rect 4019 311 4622 317
rect 4019 271 4565 311
rect 3507 265 4565 271
rect 4611 265 4622 311
rect 3507 232 3686 265
rect 4081 244 4498 265
rect 3762 173 4021 219
rect 3762 160 3808 173
rect 1262 127 1330 128
rect 446 81 457 127
rect 503 81 514 127
rect 446 60 514 81
rect 1262 81 1273 127
rect 1319 81 1330 127
rect 1262 60 1330 81
rect 2222 81 2233 127
rect 2279 81 2290 127
rect 2222 60 2290 81
rect 3038 81 3049 127
rect 3095 81 3106 127
rect 3162 114 3457 160
rect 3503 114 3808 160
rect 3975 152 4021 173
rect 4567 173 5089 219
rect 5135 173 5146 219
rect 4567 152 4613 173
rect 3038 60 3106 81
rect 3854 81 3865 127
rect 3911 81 3922 127
rect 3975 106 4273 152
rect 4319 106 4613 152
rect 4946 130 5146 173
rect 3854 60 3922 81
rect 4670 81 4681 127
rect 4727 81 4738 127
rect 4670 60 4738 81
rect 0 -60 5264 60
<< labels >>
flabel metal1 s 3556 393 5134 439 0 FreeSans 600 0 0 0 A1
port 1 nsew default input
flabel metal1 s 3415 521 4942 567 0 FreeSans 600 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 1262 127 1330 128 0 FreeSans 600 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 0 724 5264 844 0 FreeSans 600 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 117 360 1418 424 0 FreeSans 600 0 0 0 C2
port 6 nsew default input
flabel metal1 s 1464 352 1703 430 0 FreeSans 600 0 0 0 C1
port 5 nsew default input
flabel metal1 s 2083 360 3251 424 0 FreeSans 600 0 0 0 B2
port 4 nsew default input
flabel metal1 s 1789 405 2032 430 0 FreeSans 600 0 0 0 B1
port 3 nsew default input
flabel metal1 s 3507 265 4622 323 0 FreeSans 600 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 4722 354 5134 393 1 A1
port 1 nsew default input
rlabel metal1 s 4081 244 4498 265 1 A2
port 2 nsew default input
rlabel metal1 s 3507 244 3686 265 1 A2
port 2 nsew default input
rlabel metal1 s 3507 232 3686 244 1 A2
port 2 nsew default input
rlabel metal1 s 3321 313 3367 405 1 B1
port 3 nsew default input
rlabel metal1 s 1789 313 2032 405 1 B1
port 3 nsew default input
rlabel metal1 s 1789 267 3367 313 1 B1
port 3 nsew default input
rlabel metal1 s 1464 313 1524 352 1 C1
port 5 nsew default input
rlabel metal1 s 142 267 1524 313 1 C1
port 5 nsew default input
rlabel metal1 s 3415 220 3461 521 1 ZN
port 7 nsew default output
rlabel metal1 s 3415 219 3461 220 1 ZN
port 7 nsew default output
rlabel metal1 s 1126 219 1407 220 1 ZN
port 7 nsew default output
rlabel metal1 s 4567 174 5146 219 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 174 4021 219 1 ZN
port 7 nsew default output
rlabel metal1 s 3415 174 3461 219 1 ZN
port 7 nsew default output
rlabel metal1 s 38 174 3208 219 1 ZN
port 7 nsew default output
rlabel metal1 s 4567 173 5146 174 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 173 4021 174 1 ZN
port 7 nsew default output
rlabel metal1 s 3415 173 3461 174 1 ZN
port 7 nsew default output
rlabel metal1 s 1361 173 3208 174 1 ZN
port 7 nsew default output
rlabel metal1 s 38 173 1172 174 1 ZN
port 7 nsew default output
rlabel metal1 s 4946 160 5146 173 1 ZN
port 7 nsew default output
rlabel metal1 s 4567 160 4613 173 1 ZN
port 7 nsew default output
rlabel metal1 s 3975 160 4021 173 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 160 3808 173 1 ZN
port 7 nsew default output
rlabel metal1 s 3415 160 3461 173 1 ZN
port 7 nsew default output
rlabel metal1 s 3162 160 3208 173 1 ZN
port 7 nsew default output
rlabel metal1 s 4946 152 5146 160 1 ZN
port 7 nsew default output
rlabel metal1 s 4567 152 4613 160 1 ZN
port 7 nsew default output
rlabel metal1 s 3975 152 4021 160 1 ZN
port 7 nsew default output
rlabel metal1 s 3162 152 3808 160 1 ZN
port 7 nsew default output
rlabel metal1 s 4946 130 5146 152 1 ZN
port 7 nsew default output
rlabel metal1 s 3975 130 4613 152 1 ZN
port 7 nsew default output
rlabel metal1 s 3162 130 3808 152 1 ZN
port 7 nsew default output
rlabel metal1 s 3975 114 4613 130 1 ZN
port 7 nsew default output
rlabel metal1 s 3162 114 3808 130 1 ZN
port 7 nsew default output
rlabel metal1 s 3975 106 4613 114 1 ZN
port 7 nsew default output
rlabel metal1 s 1670 608 1738 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1262 608 1330 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 854 608 922 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 446 608 515 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 38 608 106 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 38 511 106 608 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4670 60 4738 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3854 60 3922 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3038 60 3106 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 2222 60 2290 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1262 60 1330 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 446 60 514 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5264 60 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5264 784
string GDS_END 1330570
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1321056
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
