magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< metal2 >>
rect 0 9169 208 9199
rect 0 9009 18 9169
rect 178 9009 208 9169
rect 0 2570 208 9009
rect 0 2410 18 2570
rect 178 2410 208 2570
rect 0 2380 208 2410
rect 358 8848 566 8880
rect 358 8688 376 8848
rect 536 8688 566 8848
rect 358 2225 566 8688
rect 358 2065 376 2225
rect 536 2065 566 2225
rect 358 2040 566 2065
rect 694 8532 902 8554
rect 694 8372 712 8532
rect 872 8372 902 8532
rect 694 1905 902 8372
rect 694 1745 712 1905
rect 872 1745 902 1905
rect 694 1700 902 1745
rect 1029 8210 1237 8235
rect 1029 8050 1049 8210
rect 1209 8050 1237 8210
rect 1029 1562 1237 8050
rect 1029 1402 1049 1562
rect 1209 1402 1237 1562
rect 1029 1360 1237 1402
rect 1369 7519 1577 7544
rect 1369 7359 1389 7519
rect 1549 7359 1577 7519
rect 1369 1228 1577 7359
rect 1369 1068 1389 1228
rect 1549 1068 1577 1228
rect 1369 1020 1577 1068
rect 1706 7198 1914 7223
rect 1706 7038 1726 7198
rect 1886 7038 1914 7198
rect 1706 855 1914 7038
rect 1706 695 1726 855
rect 1886 695 1914 855
rect 1706 681 1914 695
rect 2034 6877 2242 6902
rect 2034 6717 2054 6877
rect 2214 6717 2242 6877
rect 2034 534 2242 6717
rect 2034 374 2054 534
rect 2214 374 2242 534
rect 2034 340 2242 374
rect 2393 6551 2601 6580
rect 2393 6391 2426 6551
rect 2586 6391 2601 6551
rect 2393 195 2601 6391
rect 2393 35 2414 195
rect 2574 35 2601 195
rect 2393 0 2601 35
<< via2 >>
rect 18 9009 178 9169
rect 18 2410 178 2570
rect 376 8688 536 8848
rect 376 2065 536 2225
rect 712 8372 872 8532
rect 712 1745 872 1905
rect 1049 8050 1209 8210
rect 1049 1402 1209 1562
rect 1389 7359 1549 7519
rect 1389 1068 1549 1228
rect 1726 7038 1886 7198
rect 1726 695 1886 855
rect 2054 6717 2214 6877
rect 2054 374 2214 534
rect 2426 6391 2586 6551
rect 2414 35 2574 195
<< metal3 >>
rect 1 9169 3541 9202
rect 1 9009 18 9169
rect 178 9009 3541 9169
rect 1 8987 3541 9009
rect 358 8848 3541 8880
rect 358 8688 376 8848
rect 536 8688 3541 8848
rect 358 8665 3541 8688
rect 694 8532 3541 8559
rect 694 8372 712 8532
rect 872 8372 3541 8532
rect 694 8344 3541 8372
rect 1029 8210 3541 8237
rect 1029 8050 1049 8210
rect 1209 8050 3541 8210
rect 1029 8022 3541 8050
rect 1369 7519 3541 7545
rect 1369 7359 1389 7519
rect 1549 7359 3541 7519
rect 1369 7330 3541 7359
rect 1708 7198 3541 7223
rect 1708 7038 1726 7198
rect 1886 7038 3541 7198
rect 1708 7008 3541 7038
rect 2036 6877 3541 6902
rect 2036 6717 2054 6877
rect 2214 6717 3541 6877
rect 2036 6687 3541 6717
rect 2394 6551 3541 6579
rect 2394 6391 2426 6551
rect 2586 6391 3541 6551
rect 2394 6364 3541 6391
rect 8 2570 188 2580
rect 8 2410 18 2570
rect 178 2410 188 2570
rect 8 2400 188 2410
rect 366 2225 546 2235
rect 366 2065 376 2225
rect 536 2065 546 2225
rect 366 2055 546 2065
rect 702 1905 882 1915
rect 702 1745 712 1905
rect 872 1745 882 1905
rect 702 1735 882 1745
rect 1039 1562 1219 1572
rect 1039 1402 1049 1562
rect 1209 1402 1219 1562
rect 1039 1392 1219 1402
rect 1379 1228 1559 1238
rect 1379 1068 1389 1228
rect 1549 1068 1559 1228
rect 1379 1058 1559 1068
rect 1716 855 1896 865
rect 1716 695 1726 855
rect 1886 695 1896 855
rect 1716 685 1896 695
rect 2044 534 2224 544
rect 2044 374 2054 534
rect 2214 374 2224 534
rect 2044 364 2224 374
rect 2404 195 2584 205
rect 2404 35 2414 195
rect 2574 35 2584 195
rect 2404 25 2584 35
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1750858719
transform -1 0 98 0 1 2490
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1750858719
transform -1 0 456 0 1 2145
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1750858719
transform -1 0 792 0 1 1825
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1750858719
transform -1 0 1129 0 1 1482
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1750858719
transform -1 0 1469 0 1 1148
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1750858719
transform -1 0 1806 0 1 775
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1750858719
transform -1 0 2134 0 1 454
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1750858719
transform -1 0 2494 0 1 115
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1750858719
transform -1 0 2134 0 1 6797
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1750858719
transform -1 0 1806 0 1 7118
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1750858719
transform -1 0 1469 0 1 7439
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1750858719
transform -1 0 1129 0 1 8130
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1750858719
transform -1 0 792 0 1 8452
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1750858719
transform -1 0 456 0 1 8768
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1750858719
transform -1 0 98 0 1 9089
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1750858719
transform -1 0 2506 0 1 6471
box 0 0 1 1
<< properties >>
string GDS_END 2833688
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2831572
<< end >>
