magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< metal1 >>
rect 0 918 1120 1098
rect 487 710 533 918
rect 142 454 214 542
rect 359 443 418 542
rect 49 90 95 298
rect 497 90 543 298
rect 702 136 767 872
rect 925 710 971 918
rect 945 90 991 298
rect 0 -90 1120 90
<< obsm1 >>
rect 69 664 115 872
rect 69 618 641 664
rect 595 390 641 618
rect 273 344 641 390
rect 273 136 319 344
<< labels >>
rlabel metal1 s 142 454 214 542 6 A1
port 1 nsew default input
rlabel metal1 s 359 443 418 542 6 A2
port 2 nsew default input
rlabel metal1 s 702 136 767 872 6 Z
port 3 nsew default output
rlabel metal1 s 925 710 971 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 487 710 533 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 918 1120 1098 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s -86 453 1206 1094 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 1206 453 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -90 1120 90 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 298 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 269876
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 266240
<< end >>
