magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3520 1660
<< nmos >>
rect 190 210 250 380
rect 540 210 600 380
rect 710 210 770 380
rect 1060 210 1120 380
rect 1220 210 1280 380
rect 1390 210 1450 380
rect 1500 210 1560 380
rect 1670 210 1730 380
rect 1780 210 1840 380
rect 1950 210 2010 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2580 210 2640 380
rect 2750 210 2810 380
rect 3100 210 3160 380
rect 3270 210 3330 380
<< pmos >>
rect 190 1110 250 1450
rect 510 1110 570 1450
rect 620 1110 680 1450
rect 1060 1110 1120 1450
rect 1220 1110 1280 1450
rect 1390 1110 1450 1450
rect 1500 1110 1560 1450
rect 1670 1110 1730 1450
rect 1780 1110 1840 1450
rect 1950 1110 2010 1450
rect 2060 1110 2120 1450
rect 2230 1110 2290 1450
rect 2670 1110 2730 1450
rect 2780 1110 2840 1450
rect 3100 1110 3160 1450
rect 3270 1110 3330 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 440 318 540 380
rect 440 272 462 318
rect 508 272 540 318
rect 440 210 540 272
rect 600 318 710 380
rect 600 272 632 318
rect 678 272 710 318
rect 600 210 710 272
rect 770 318 870 380
rect 770 272 802 318
rect 848 272 870 318
rect 770 210 870 272
rect 960 318 1060 380
rect 960 272 982 318
rect 1028 272 1060 318
rect 960 210 1060 272
rect 1120 210 1220 380
rect 1280 318 1390 380
rect 1280 272 1312 318
rect 1358 272 1390 318
rect 1280 210 1390 272
rect 1450 210 1500 380
rect 1560 278 1670 380
rect 1560 232 1592 278
rect 1638 232 1670 278
rect 1560 210 1670 232
rect 1730 210 1780 380
rect 1840 318 1950 380
rect 1840 272 1872 318
rect 1918 272 1950 318
rect 1840 210 1950 272
rect 2010 210 2060 380
rect 2120 318 2230 380
rect 2120 272 2152 318
rect 2198 272 2230 318
rect 2120 210 2230 272
rect 2290 318 2390 380
rect 2290 272 2322 318
rect 2368 272 2390 318
rect 2290 210 2390 272
rect 2480 318 2580 380
rect 2480 272 2502 318
rect 2548 272 2580 318
rect 2480 210 2580 272
rect 2640 318 2750 380
rect 2640 272 2672 318
rect 2718 272 2750 318
rect 2640 210 2750 272
rect 2810 318 2910 380
rect 2810 272 2842 318
rect 2888 272 2910 318
rect 2810 210 2910 272
rect 3000 318 3100 380
rect 3000 272 3022 318
rect 3068 272 3100 318
rect 3000 210 3100 272
rect 3160 318 3270 380
rect 3160 272 3192 318
rect 3238 272 3270 318
rect 3160 210 3270 272
rect 3330 318 3430 380
rect 3330 272 3362 318
rect 3408 272 3430 318
rect 3330 210 3430 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 350 1450
rect 250 1163 282 1397
rect 328 1163 350 1397
rect 250 1110 350 1163
rect 410 1397 510 1450
rect 410 1163 432 1397
rect 478 1163 510 1397
rect 410 1110 510 1163
rect 570 1110 620 1450
rect 680 1397 780 1450
rect 680 1163 712 1397
rect 758 1163 780 1397
rect 680 1110 780 1163
rect 960 1397 1060 1450
rect 960 1163 982 1397
rect 1028 1163 1060 1397
rect 960 1110 1060 1163
rect 1120 1110 1220 1450
rect 1280 1397 1390 1450
rect 1280 1163 1312 1397
rect 1358 1163 1390 1397
rect 1280 1110 1390 1163
rect 1450 1110 1500 1450
rect 1560 1397 1670 1450
rect 1560 1163 1592 1397
rect 1638 1163 1670 1397
rect 1560 1110 1670 1163
rect 1730 1110 1780 1450
rect 1840 1425 1950 1450
rect 1840 1285 1872 1425
rect 1918 1285 1950 1425
rect 1840 1110 1950 1285
rect 2010 1110 2060 1450
rect 2120 1425 2230 1450
rect 2120 1285 2152 1425
rect 2198 1285 2230 1425
rect 2120 1110 2230 1285
rect 2290 1397 2390 1450
rect 2290 1163 2322 1397
rect 2368 1163 2390 1397
rect 2290 1110 2390 1163
rect 2570 1397 2670 1450
rect 2570 1163 2592 1397
rect 2638 1163 2670 1397
rect 2570 1110 2670 1163
rect 2730 1110 2780 1450
rect 2840 1397 2940 1450
rect 2840 1163 2872 1397
rect 2918 1163 2940 1397
rect 2840 1110 2940 1163
rect 3000 1397 3100 1450
rect 3000 1163 3022 1397
rect 3068 1163 3100 1397
rect 3000 1110 3100 1163
rect 3160 1397 3270 1450
rect 3160 1163 3192 1397
rect 3238 1163 3270 1397
rect 3160 1110 3270 1163
rect 3330 1397 3430 1450
rect 3330 1163 3362 1397
rect 3408 1163 3430 1397
rect 3330 1110 3430 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 462 272 508 318
rect 632 272 678 318
rect 802 272 848 318
rect 982 272 1028 318
rect 1312 272 1358 318
rect 1592 232 1638 278
rect 1872 272 1918 318
rect 2152 272 2198 318
rect 2322 272 2368 318
rect 2502 272 2548 318
rect 2672 272 2718 318
rect 2842 272 2888 318
rect 3022 272 3068 318
rect 3192 272 3238 318
rect 3362 272 3408 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 432 1163 478 1397
rect 712 1163 758 1397
rect 982 1163 1028 1397
rect 1312 1163 1358 1397
rect 1592 1163 1638 1397
rect 1872 1285 1918 1425
rect 2152 1285 2198 1425
rect 2322 1163 2368 1397
rect 2592 1163 2638 1397
rect 2872 1163 2918 1397
rect 3022 1163 3068 1397
rect 3192 1163 3238 1397
rect 3362 1163 3408 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 560 118 710 140
rect 560 72 612 118
rect 658 72 710 118
rect 560 50 710 72
rect 810 118 960 140
rect 810 72 862 118
rect 908 72 960 118
rect 810 50 960 72
rect 1060 118 1210 140
rect 1060 72 1112 118
rect 1158 72 1210 118
rect 1060 50 1210 72
rect 1310 118 1460 140
rect 1310 72 1362 118
rect 1408 72 1460 118
rect 1310 50 1460 72
rect 1560 118 1710 140
rect 1560 72 1612 118
rect 1658 72 1710 118
rect 1560 50 1710 72
rect 1810 118 1960 140
rect 1810 72 1862 118
rect 1908 72 1960 118
rect 1810 50 1960 72
rect 2060 118 2210 140
rect 2060 72 2112 118
rect 2158 72 2210 118
rect 2060 50 2210 72
rect 2310 118 2460 140
rect 2310 72 2362 118
rect 2408 72 2460 118
rect 2310 50 2460 72
rect 2560 118 2710 140
rect 2560 72 2612 118
rect 2658 72 2710 118
rect 2560 50 2710 72
rect 2810 118 2960 140
rect 2810 72 2862 118
rect 2908 72 2960 118
rect 2810 50 2960 72
rect 3060 118 3210 140
rect 3060 72 3112 118
rect 3158 72 3210 118
rect 3060 50 3210 72
rect 3310 118 3460 140
rect 3310 72 3362 118
rect 3408 72 3460 118
rect 3310 50 3460 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
rect 980 1588 1130 1610
rect 980 1542 1032 1588
rect 1078 1542 1130 1588
rect 980 1520 1130 1542
rect 1210 1588 1360 1610
rect 1210 1542 1262 1588
rect 1308 1542 1360 1588
rect 1210 1520 1360 1542
rect 1440 1588 1590 1610
rect 1440 1542 1492 1588
rect 1538 1542 1590 1588
rect 1440 1520 1590 1542
rect 1670 1588 1820 1610
rect 1670 1542 1722 1588
rect 1768 1542 1820 1588
rect 1670 1520 1820 1542
rect 1900 1588 2050 1610
rect 1900 1542 1952 1588
rect 1998 1542 2050 1588
rect 1900 1520 2050 1542
rect 2130 1588 2280 1610
rect 2130 1542 2182 1588
rect 2228 1542 2280 1588
rect 2130 1520 2280 1542
rect 2360 1588 2510 1610
rect 2360 1542 2412 1588
rect 2458 1542 2510 1588
rect 2360 1520 2510 1542
rect 2590 1588 2740 1610
rect 2590 1542 2642 1588
rect 2688 1542 2740 1588
rect 2590 1520 2740 1542
rect 2820 1588 2970 1610
rect 2820 1542 2872 1588
rect 2918 1542 2970 1588
rect 2820 1520 2970 1542
rect 3050 1588 3200 1610
rect 3050 1542 3102 1588
rect 3148 1542 3200 1588
rect 3050 1520 3200 1542
rect 3280 1588 3430 1610
rect 3280 1542 3332 1588
rect 3378 1542 3430 1588
rect 3280 1520 3430 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 612 72 658 118
rect 862 72 908 118
rect 1112 72 1158 118
rect 1362 72 1408 118
rect 1612 72 1658 118
rect 1862 72 1908 118
rect 2112 72 2158 118
rect 2362 72 2408 118
rect 2612 72 2658 118
rect 2862 72 2908 118
rect 3112 72 3158 118
rect 3362 72 3408 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
rect 1032 1542 1078 1588
rect 1262 1542 1308 1588
rect 1492 1542 1538 1588
rect 1722 1542 1768 1588
rect 1952 1542 1998 1588
rect 2182 1542 2228 1588
rect 2412 1542 2458 1588
rect 2642 1542 2688 1588
rect 2872 1542 2918 1588
rect 3102 1542 3148 1588
rect 3332 1542 3378 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 510 1450 570 1500
rect 620 1450 680 1500
rect 1060 1450 1120 1500
rect 1220 1450 1280 1500
rect 1390 1450 1450 1500
rect 1500 1450 1560 1500
rect 1670 1450 1730 1500
rect 1780 1450 1840 1500
rect 1950 1450 2010 1500
rect 2060 1450 2120 1500
rect 2230 1450 2290 1500
rect 2670 1450 2730 1500
rect 2780 1450 2840 1500
rect 3100 1450 3160 1500
rect 3270 1450 3330 1500
rect 190 1060 250 1110
rect 120 1038 250 1060
rect 120 992 142 1038
rect 188 992 250 1038
rect 120 970 250 992
rect 190 380 250 970
rect 510 800 570 1110
rect 620 1060 680 1110
rect 620 1000 770 1060
rect 710 930 770 1000
rect 710 903 880 930
rect 710 857 797 903
rect 843 857 880 903
rect 710 830 880 857
rect 510 773 630 800
rect 510 727 557 773
rect 603 727 630 773
rect 510 700 630 727
rect 510 650 570 700
rect 510 610 600 650
rect 540 380 600 610
rect 710 380 770 830
rect 1060 800 1120 1110
rect 1220 930 1280 1110
rect 1220 903 1320 930
rect 1220 857 1247 903
rect 1293 857 1320 903
rect 1220 830 1320 857
rect 1060 773 1180 800
rect 1060 727 1107 773
rect 1153 727 1180 773
rect 1060 700 1180 727
rect 1060 380 1120 700
rect 1390 660 1450 1110
rect 1500 1060 1560 1110
rect 1670 1060 1730 1110
rect 1500 1033 1730 1060
rect 1500 990 1537 1033
rect 1510 987 1537 990
rect 1583 990 1730 1033
rect 1583 987 1610 990
rect 1510 940 1610 987
rect 1780 660 1840 1110
rect 1950 930 2010 1110
rect 1910 903 2010 930
rect 1910 857 1937 903
rect 1983 857 2010 903
rect 1910 830 2010 857
rect 2060 800 2120 1110
rect 2230 930 2290 1110
rect 2670 1060 2730 1110
rect 2550 1000 2730 1060
rect 2230 903 2330 930
rect 2230 857 2257 903
rect 2303 857 2330 903
rect 2230 830 2330 857
rect 2050 773 2150 800
rect 2050 727 2077 773
rect 2123 727 2150 773
rect 2050 700 2150 727
rect 1910 660 2010 670
rect 1220 643 2010 660
rect 1220 600 1937 643
rect 1220 380 1280 600
rect 1910 597 1937 600
rect 1983 597 2010 643
rect 1910 570 2010 597
rect 1350 513 1450 540
rect 1510 520 1610 540
rect 1350 467 1377 513
rect 1423 467 1450 513
rect 1350 440 1450 467
rect 1390 380 1450 440
rect 1500 513 1730 520
rect 1500 467 1537 513
rect 1583 467 1730 513
rect 1500 440 1730 467
rect 1500 380 1560 440
rect 1670 380 1730 440
rect 1780 503 1880 530
rect 1780 457 1807 503
rect 1853 457 1880 503
rect 1780 430 1880 457
rect 1780 380 1840 430
rect 1950 380 2010 570
rect 2060 380 2120 700
rect 2230 380 2290 830
rect 2550 530 2610 1000
rect 2780 650 2840 1110
rect 3100 670 3160 1110
rect 3270 930 3330 1110
rect 3210 903 3330 930
rect 3210 857 3237 903
rect 3283 857 3330 903
rect 3210 830 3330 857
rect 2470 503 2610 530
rect 2470 457 2507 503
rect 2553 470 2610 503
rect 2750 610 2840 650
rect 3040 643 3160 670
rect 2750 530 2810 610
rect 3040 597 3087 643
rect 3133 597 3160 643
rect 3040 570 3160 597
rect 2750 503 2870 530
rect 2553 457 2640 470
rect 2470 430 2640 457
rect 2580 380 2640 430
rect 2750 457 2797 503
rect 2843 457 2870 503
rect 2750 430 2870 457
rect 2750 380 2810 430
rect 3100 380 3160 570
rect 3270 380 3330 830
rect 190 160 250 210
rect 540 160 600 210
rect 710 160 770 210
rect 1060 160 1120 210
rect 1220 160 1280 210
rect 1390 160 1450 210
rect 1500 160 1560 210
rect 1670 160 1730 210
rect 1780 160 1840 210
rect 1950 160 2010 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2580 160 2640 210
rect 2750 160 2810 210
rect 3100 160 3160 210
rect 3270 160 3330 210
<< polycontact >>
rect 142 992 188 1038
rect 797 857 843 903
rect 557 727 603 773
rect 1247 857 1293 903
rect 1107 727 1153 773
rect 1537 987 1583 1033
rect 1937 857 1983 903
rect 2257 857 2303 903
rect 2077 727 2123 773
rect 1937 597 1983 643
rect 1377 467 1423 513
rect 1537 467 1583 513
rect 1807 457 1853 503
rect 3237 857 3283 903
rect 2507 457 2553 503
rect 3087 597 3133 643
rect 2797 457 2843 503
<< metal1 >>
rect 0 1588 3520 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1032 1588
rect 1078 1542 1262 1588
rect 1308 1542 1492 1588
rect 1538 1542 1722 1588
rect 1768 1542 1952 1588
rect 1998 1542 2182 1588
rect 2228 1542 2412 1588
rect 2458 1542 2642 1588
rect 2688 1542 2872 1588
rect 2918 1542 3102 1588
rect 3148 1542 3332 1588
rect 3378 1542 3520 1588
rect 0 1520 3520 1542
rect 110 1397 160 1520
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1110 160 1163
rect 280 1397 330 1450
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 110 1038 210 1040
rect 110 1036 142 1038
rect 110 984 134 1036
rect 188 992 210 1038
rect 186 984 210 992
rect 110 980 210 984
rect 280 520 330 1163
rect 430 1397 480 1450
rect 430 1163 432 1397
rect 478 1163 480 1397
rect 430 570 480 1163
rect 710 1397 760 1520
rect 710 1163 712 1397
rect 758 1163 760 1397
rect 710 1110 760 1163
rect 980 1397 1030 1520
rect 980 1163 982 1397
rect 1028 1163 1030 1397
rect 980 1110 1030 1163
rect 1310 1397 1360 1450
rect 1310 1163 1312 1397
rect 1358 1163 1360 1397
rect 1310 1060 1360 1163
rect 1590 1397 1640 1520
rect 1590 1163 1592 1397
rect 1638 1163 1640 1397
rect 1870 1425 1920 1450
rect 1870 1285 1872 1425
rect 1918 1285 1920 1425
rect 1870 1260 1920 1285
rect 2150 1425 2200 1520
rect 2150 1285 2152 1425
rect 2198 1285 2200 1425
rect 2150 1260 2200 1285
rect 2320 1397 2370 1450
rect 1590 1110 1640 1163
rect 1690 1210 1920 1260
rect 980 1010 1360 1060
rect 1510 1033 1610 1040
rect 980 910 1030 1010
rect 1510 987 1537 1033
rect 1583 987 1610 1033
rect 1510 980 1610 987
rect 770 903 1030 910
rect 770 857 797 903
rect 843 857 1030 903
rect 770 850 1030 857
rect 1220 906 1450 910
rect 1220 903 1374 906
rect 1220 857 1247 903
rect 1293 857 1374 903
rect 1220 854 1374 857
rect 1426 854 1450 906
rect 1220 850 1450 854
rect 530 776 630 780
rect 530 724 554 776
rect 606 724 630 776
rect 530 720 630 724
rect 430 520 680 570
rect 790 520 840 530
rect 980 520 1030 850
rect 1080 776 1180 780
rect 1080 724 1104 776
rect 1156 724 1180 776
rect 1080 720 1180 724
rect 1370 520 1430 850
rect 1530 520 1590 980
rect 1690 760 1740 1210
rect 2320 1163 2322 1397
rect 2368 1163 2370 1397
rect 2040 1036 2140 1040
rect 2040 984 2064 1036
rect 2116 984 2140 1036
rect 2040 980 2140 984
rect 2320 1020 2370 1163
rect 2590 1397 2640 1520
rect 2590 1163 2592 1397
rect 2638 1163 2640 1397
rect 2590 1110 2640 1163
rect 2870 1397 2920 1450
rect 2870 1163 2872 1397
rect 2918 1163 2920 1397
rect 2500 1040 2560 1060
rect 2870 1040 2920 1163
rect 3020 1397 3070 1450
rect 3020 1163 3022 1397
rect 3068 1163 3070 1397
rect 2500 1036 2950 1040
rect 1680 710 1740 760
rect 1800 906 2010 910
rect 1800 854 1934 906
rect 1986 854 2010 906
rect 1800 850 2010 854
rect 260 516 360 520
rect 260 464 284 516
rect 336 464 360 516
rect 260 460 360 464
rect 600 516 870 520
rect 600 464 794 516
rect 846 464 870 516
rect 980 470 1180 520
rect 600 460 870 464
rect 280 450 340 460
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 450
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 460 318 510 380
rect 460 272 462 318
rect 508 272 510 318
rect 460 140 510 272
rect 630 318 680 460
rect 790 450 840 460
rect 1100 380 1180 470
rect 1350 513 1450 520
rect 1350 467 1377 513
rect 1423 467 1450 513
rect 1350 460 1450 467
rect 1510 516 1610 520
rect 1510 464 1534 516
rect 1586 464 1610 516
rect 1510 460 1610 464
rect 1680 390 1730 710
rect 1800 510 1860 850
rect 2060 780 2120 980
rect 2320 970 2430 1020
rect 2230 906 2330 910
rect 2230 854 2254 906
rect 2306 854 2330 906
rect 2230 850 2330 854
rect 2380 780 2430 970
rect 2500 984 2504 1036
rect 2556 984 2874 1036
rect 2926 984 2950 1036
rect 2500 980 2950 984
rect 2500 960 2560 980
rect 2050 776 2150 780
rect 2050 724 2074 776
rect 2126 724 2150 776
rect 2050 720 2150 724
rect 2320 730 2430 780
rect 1910 646 2010 650
rect 1910 594 1934 646
rect 1986 594 2010 646
rect 1910 590 2010 594
rect 2320 646 2380 730
rect 2870 650 2920 980
rect 3020 910 3070 1163
rect 3190 1397 3240 1520
rect 3190 1163 3192 1397
rect 3238 1163 3240 1397
rect 3190 1110 3240 1163
rect 3360 1397 3410 1450
rect 3360 1163 3362 1397
rect 3408 1163 3410 1397
rect 3360 1050 3410 1163
rect 3360 1036 3460 1050
rect 3360 984 3384 1036
rect 3436 984 3460 1036
rect 3360 980 3460 984
rect 3360 970 3450 980
rect 3020 906 3310 910
rect 3020 854 3234 906
rect 3286 854 3310 906
rect 3020 850 3310 854
rect 2320 594 2324 646
rect 2376 594 2380 646
rect 2320 570 2380 594
rect 2670 646 3160 650
rect 2670 594 3084 646
rect 3136 594 3160 646
rect 2670 590 3160 594
rect 1780 503 1880 510
rect 1780 457 1807 503
rect 1853 457 1880 503
rect 1780 450 1880 457
rect 1680 386 1950 390
rect 630 272 632 318
rect 678 272 680 318
rect 630 210 680 272
rect 800 318 850 380
rect 800 272 802 318
rect 848 272 850 318
rect 800 140 850 272
rect 980 318 1030 380
rect 1100 330 1360 380
rect 1680 340 1874 386
rect 980 272 982 318
rect 1028 272 1030 318
rect 980 140 1030 272
rect 1310 318 1360 330
rect 1310 272 1312 318
rect 1358 272 1360 318
rect 1870 334 1874 340
rect 1926 334 1950 386
rect 1870 330 1950 334
rect 1870 318 1920 330
rect 1310 210 1360 272
rect 1590 278 1640 300
rect 1590 232 1592 278
rect 1638 232 1640 278
rect 1590 140 1640 232
rect 1870 272 1872 318
rect 1918 272 1920 318
rect 1870 210 1920 272
rect 2150 318 2200 380
rect 2150 272 2152 318
rect 2198 272 2200 318
rect 2150 140 2200 272
rect 2320 318 2370 570
rect 2480 506 2580 510
rect 2480 454 2504 506
rect 2556 454 2580 506
rect 2480 450 2580 454
rect 2320 272 2322 318
rect 2368 272 2370 318
rect 2320 210 2370 272
rect 2500 318 2550 380
rect 2500 272 2502 318
rect 2548 272 2550 318
rect 2500 140 2550 272
rect 2670 318 2720 590
rect 2770 506 2870 510
rect 2770 454 2794 506
rect 2846 454 2870 506
rect 3240 480 3290 850
rect 2770 450 2870 454
rect 3020 430 3290 480
rect 2670 272 2672 318
rect 2718 272 2720 318
rect 2670 210 2720 272
rect 2840 318 2890 380
rect 2840 272 2842 318
rect 2888 272 2890 318
rect 2840 140 2890 272
rect 3020 318 3070 430
rect 3020 272 3022 318
rect 3068 272 3070 318
rect 3020 210 3070 272
rect 3190 318 3240 380
rect 3190 272 3192 318
rect 3238 272 3240 318
rect 3190 140 3240 272
rect 3360 318 3410 970
rect 3360 272 3362 318
rect 3408 272 3410 318
rect 3360 210 3410 272
rect 0 118 3520 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 612 118
rect 658 72 862 118
rect 908 72 1112 118
rect 1158 72 1362 118
rect 1408 72 1612 118
rect 1658 72 1862 118
rect 1908 72 2112 118
rect 2158 72 2362 118
rect 2408 72 2612 118
rect 2658 72 2862 118
rect 2908 72 3112 118
rect 3158 72 3362 118
rect 3408 72 3520 118
rect 0 0 3520 72
<< via1 >>
rect 134 992 142 1036
rect 142 992 186 1036
rect 134 984 186 992
rect 1374 854 1426 906
rect 554 773 606 776
rect 554 727 557 773
rect 557 727 603 773
rect 603 727 606 773
rect 554 724 606 727
rect 1104 773 1156 776
rect 1104 727 1107 773
rect 1107 727 1153 773
rect 1153 727 1156 773
rect 1104 724 1156 727
rect 2064 984 2116 1036
rect 1934 903 1986 906
rect 1934 857 1937 903
rect 1937 857 1983 903
rect 1983 857 1986 903
rect 1934 854 1986 857
rect 284 464 336 516
rect 794 464 846 516
rect 1534 513 1586 516
rect 1534 467 1537 513
rect 1537 467 1583 513
rect 1583 467 1586 513
rect 1534 464 1586 467
rect 2254 903 2306 906
rect 2254 857 2257 903
rect 2257 857 2303 903
rect 2303 857 2306 903
rect 2254 854 2306 857
rect 2504 984 2556 1036
rect 2874 984 2926 1036
rect 2074 773 2126 776
rect 2074 727 2077 773
rect 2077 727 2123 773
rect 2123 727 2126 773
rect 2074 724 2126 727
rect 1934 643 1986 646
rect 1934 597 1937 643
rect 1937 597 1983 643
rect 1983 597 1986 643
rect 1934 594 1986 597
rect 3384 984 3436 1036
rect 3234 903 3286 906
rect 3234 857 3237 903
rect 3237 857 3283 903
rect 3283 857 3286 903
rect 3234 854 3286 857
rect 2324 594 2376 646
rect 3084 643 3136 646
rect 3084 597 3087 643
rect 3087 597 3133 643
rect 3133 597 3136 643
rect 3084 594 3136 597
rect 1874 334 1926 386
rect 2504 503 2556 506
rect 2504 457 2507 503
rect 2507 457 2553 503
rect 2553 457 2556 503
rect 2504 454 2556 457
rect 2794 503 2846 506
rect 2794 457 2797 503
rect 2797 457 2843 503
rect 2843 457 2846 503
rect 2794 454 2846 457
<< metal2 >>
rect 110 1036 210 1050
rect 2050 1040 2130 1050
rect 2490 1040 2570 1050
rect 110 984 134 1036
rect 186 984 210 1036
rect 110 970 210 984
rect 2040 1036 2580 1040
rect 2040 984 2064 1036
rect 2116 984 2504 1036
rect 2556 984 2580 1036
rect 2040 980 2580 984
rect 2850 1036 2950 1050
rect 3370 1040 3450 1050
rect 2850 984 2874 1036
rect 2926 984 2950 1036
rect 2050 970 2130 980
rect 2490 970 2570 980
rect 2850 970 2950 984
rect 3360 1036 3460 1040
rect 3360 984 3384 1036
rect 3436 984 3460 1036
rect 3360 980 3460 984
rect 3370 970 3450 980
rect 1350 910 1440 920
rect 1910 910 2010 920
rect 2240 910 2320 920
rect 3220 910 3300 920
rect 1350 906 2330 910
rect 1350 854 1374 906
rect 1426 854 1934 906
rect 1986 854 2254 906
rect 2306 854 2330 906
rect 1350 850 2330 854
rect 3210 906 3310 910
rect 3210 854 3234 906
rect 3286 854 3310 906
rect 3210 850 3310 854
rect 1350 840 1440 850
rect 1910 840 2010 850
rect 2240 840 2320 850
rect 3220 840 3300 850
rect 530 776 630 790
rect 530 724 554 776
rect 606 724 630 776
rect 530 710 630 724
rect 1080 776 1180 790
rect 2060 780 2140 790
rect 1080 724 1104 776
rect 1156 724 1180 776
rect 1080 710 1180 724
rect 2050 776 2150 780
rect 2050 724 2074 776
rect 2126 724 2150 776
rect 2050 720 2150 724
rect 2060 710 2140 720
rect 260 520 360 530
rect 550 520 610 710
rect 1920 650 2000 660
rect 2310 650 2390 660
rect 3070 650 3150 660
rect 1910 646 2410 650
rect 1910 594 1934 646
rect 1986 594 2324 646
rect 2376 594 2410 646
rect 1910 590 2410 594
rect 3000 646 3160 650
rect 3000 594 3084 646
rect 3136 594 3160 646
rect 3000 590 3160 594
rect 1920 580 2000 590
rect 2310 580 2390 590
rect 3070 580 3150 590
rect 260 516 610 520
rect 260 464 284 516
rect 336 464 610 516
rect 260 460 610 464
rect 260 450 360 460
rect 550 260 610 460
rect 770 520 870 530
rect 1520 520 1600 530
rect 770 516 1610 520
rect 770 464 794 516
rect 846 464 1534 516
rect 1586 464 1610 516
rect 770 460 1610 464
rect 2480 506 2580 520
rect 770 450 870 460
rect 1520 450 1600 460
rect 2480 454 2504 506
rect 2556 454 2580 506
rect 2480 440 2580 454
rect 2750 506 2870 520
rect 2750 454 2794 506
rect 2846 454 2870 506
rect 2750 440 2870 454
rect 1860 390 1940 400
rect 2480 390 2560 440
rect 1850 386 2560 390
rect 1850 334 1874 386
rect 1926 334 2560 386
rect 1850 330 2560 334
rect 1860 320 1940 330
rect 2750 260 2810 440
rect 550 200 2810 260
<< labels >>
rlabel via1 s 1104 724 1156 776 4 D
port 1 nsew signal input
rlabel via1 s 3384 984 3436 1036 4 Q
port 2 nsew signal output
rlabel via1 s 3234 854 3286 906 4 QN
port 3 nsew signal output
rlabel via1 s 2254 854 2306 906 4 CLK
port 4 nsew clock input
rlabel via1 s 134 984 186 1036 4 RN
port 5 nsew signal input
rlabel metal1 s 110 1110 160 1660 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 710 1110 760 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 980 1110 1030 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1590 1110 1640 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 1260 2200 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2590 1110 2640 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3190 1110 3240 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3520 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 460 0 510 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 800 0 850 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 980 0 1030 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1590 0 1640 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2150 0 2200 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2500 0 2550 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2840 0 2890 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3190 0 3240 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3520 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel via1 s 1934 854 1986 906 1 CLK
port 4 nsew clock input
rlabel via1 s 1374 854 1426 906 1 CLK
port 4 nsew clock input
rlabel metal2 s 1350 840 1440 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 1910 840 2010 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 2240 840 2320 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 1350 850 2330 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1370 460 1430 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1350 460 1450 520 1 CLK
port 4 nsew clock input
rlabel metal1 s 1220 850 1450 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1800 450 1860 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1780 450 1880 510 1 CLK
port 4 nsew clock input
rlabel metal1 s 1800 850 2010 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 2230 850 2330 910 1 CLK
port 4 nsew clock input
rlabel metal2 s 1080 710 1180 790 1 D
port 1 nsew signal input
rlabel metal1 s 1080 720 1180 780 1 D
port 1 nsew signal input
rlabel metal2 s 3370 970 3450 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3360 980 3460 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 3360 210 3410 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 3360 970 3450 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 3360 980 3460 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3220 840 3300 920 1 QN
port 3 nsew signal output
rlabel metal2 s 3210 850 3310 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3020 210 3070 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3020 850 3070 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 3020 430 3290 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3240 430 3290 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3020 850 3310 910 1 QN
port 3 nsew signal output
rlabel metal2 s 110 970 210 1050 1 RN
port 5 nsew signal input
rlabel metal1 s 110 980 210 1040 1 RN
port 5 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 3520 1660
string GDS_END 238976
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 212524
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
