magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 3670 870
<< pwell >>
rect -86 -86 3670 352
<< mvnmos >>
rect 124 156 244 229
rect 348 156 468 229
rect 592 156 712 229
rect 821 156 941 229
rect 1081 156 1201 232
rect 1537 156 1657 229
rect 1781 156 1901 229
rect 2177 156 2297 229
rect 2401 156 2521 229
rect 2625 156 2745 229
rect 2849 156 2969 229
rect 3073 156 3193 229
rect 3297 156 3417 229
<< mvpmos >>
rect 124 515 224 628
rect 396 515 496 628
rect 628 515 728 628
rect 841 515 941 628
rect 1081 472 1181 628
rect 1525 515 1625 628
rect 1801 515 1901 628
rect 2197 515 2297 628
rect 2421 515 2521 628
rect 2625 515 2725 628
rect 2829 515 2929 628
rect 3073 515 3173 628
rect 3297 515 3397 628
<< mvndiff >>
rect 1001 229 1081 232
rect 36 215 124 229
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 229
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 215 592 229
rect 468 169 497 215
rect 543 169 592 215
rect 468 156 592 169
rect 712 215 821 229
rect 712 169 746 215
rect 792 169 821 215
rect 712 156 821 169
rect 941 215 1081 229
rect 941 169 970 215
rect 1016 169 1081 215
rect 941 156 1081 169
rect 1201 215 1289 232
rect 1201 169 1230 215
rect 1276 169 1289 215
rect 1201 156 1289 169
rect 1392 215 1537 229
rect 1392 169 1405 215
rect 1451 169 1537 215
rect 1392 156 1537 169
rect 1657 215 1781 229
rect 1657 169 1706 215
rect 1752 169 1781 215
rect 1657 156 1781 169
rect 1901 215 1989 229
rect 1901 169 1930 215
rect 1976 169 1989 215
rect 1901 156 1989 169
rect 2089 216 2177 229
rect 2089 170 2102 216
rect 2148 170 2177 216
rect 2089 156 2177 170
rect 2297 216 2401 229
rect 2297 170 2326 216
rect 2372 170 2401 216
rect 2297 156 2401 170
rect 2521 216 2625 229
rect 2521 170 2550 216
rect 2596 170 2625 216
rect 2521 156 2625 170
rect 2745 216 2849 229
rect 2745 170 2774 216
rect 2820 170 2849 216
rect 2745 156 2849 170
rect 2969 216 3073 229
rect 2969 170 2998 216
rect 3044 170 3073 216
rect 2969 156 3073 170
rect 3193 216 3297 229
rect 3193 170 3222 216
rect 3268 170 3297 216
rect 3193 156 3297 170
rect 3417 216 3505 229
rect 3417 170 3446 216
rect 3492 170 3505 216
rect 3417 156 3505 170
<< mvpdiff >>
rect 36 594 124 628
rect 36 548 49 594
rect 95 548 124 594
rect 36 515 124 548
rect 224 594 396 628
rect 224 548 253 594
rect 299 548 396 594
rect 224 515 396 548
rect 496 594 628 628
rect 496 548 538 594
rect 584 548 628 594
rect 496 515 628 548
rect 728 574 841 628
rect 728 528 757 574
rect 803 528 841 574
rect 728 515 841 528
rect 941 615 1081 628
rect 941 569 980 615
rect 1026 569 1081 615
rect 941 515 1081 569
rect 1001 472 1081 515
rect 1181 571 1269 628
rect 1181 525 1210 571
rect 1256 525 1269 571
rect 1181 472 1269 525
rect 1395 590 1525 628
rect 1395 544 1408 590
rect 1454 544 1525 590
rect 1395 515 1525 544
rect 1625 590 1801 628
rect 1625 544 1694 590
rect 1740 544 1801 590
rect 1625 515 1801 544
rect 1901 590 1989 628
rect 1901 544 1930 590
rect 1976 544 1989 590
rect 1901 515 1989 544
rect 2109 574 2197 628
rect 2109 528 2122 574
rect 2168 528 2197 574
rect 2109 515 2197 528
rect 2297 615 2421 628
rect 2297 569 2346 615
rect 2392 569 2421 615
rect 2297 515 2421 569
rect 2521 574 2625 628
rect 2521 528 2550 574
rect 2596 528 2625 574
rect 2521 515 2625 528
rect 2725 574 2829 628
rect 2725 528 2754 574
rect 2800 528 2829 574
rect 2725 515 2829 528
rect 2929 609 3073 628
rect 2929 563 2981 609
rect 3027 563 3073 609
rect 2929 515 3073 563
rect 3173 609 3297 628
rect 3173 563 3202 609
rect 3248 563 3297 609
rect 3173 515 3297 563
rect 3397 609 3485 628
rect 3397 563 3426 609
rect 3472 563 3485 609
rect 3397 515 3485 563
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 497 169 543 215
rect 746 169 792 215
rect 970 169 1016 215
rect 1230 169 1276 215
rect 1405 169 1451 215
rect 1706 169 1752 215
rect 1930 169 1976 215
rect 2102 170 2148 216
rect 2326 170 2372 216
rect 2550 170 2596 216
rect 2774 170 2820 216
rect 2998 170 3044 216
rect 3222 170 3268 216
rect 3446 170 3492 216
<< mvpdiffc >>
rect 49 548 95 594
rect 253 548 299 594
rect 538 548 584 594
rect 757 528 803 574
rect 980 569 1026 615
rect 1210 525 1256 571
rect 1408 544 1454 590
rect 1694 544 1740 590
rect 1930 544 1976 590
rect 2122 528 2168 574
rect 2346 569 2392 615
rect 2550 528 2596 574
rect 2754 528 2800 574
rect 2981 563 3027 609
rect 3202 563 3248 609
rect 3426 563 3472 609
<< polysilicon >>
rect 628 720 2725 760
rect 124 628 224 672
rect 396 628 496 672
rect 628 628 728 720
rect 841 628 941 672
rect 1081 628 1181 672
rect 1525 628 1625 672
rect 1801 628 1901 672
rect 2197 628 2297 672
rect 2421 628 2521 672
rect 2625 628 2725 720
rect 2829 720 3397 760
rect 2829 628 2929 720
rect 3073 628 3173 672
rect 3297 628 3397 720
rect 124 420 224 515
rect 396 482 496 515
rect 396 436 437 482
rect 483 436 496 482
rect 396 423 496 436
rect 124 394 244 420
rect 628 409 728 515
rect 841 415 941 515
rect 124 348 141 394
rect 187 348 244 394
rect 544 369 728 409
rect 821 394 941 415
rect 544 361 592 369
rect 124 229 244 348
rect 348 321 592 361
rect 821 348 865 394
rect 911 348 941 394
rect 348 229 468 321
rect 640 308 712 321
rect 640 273 653 308
rect 592 262 653 273
rect 699 262 712 308
rect 592 229 712 262
rect 821 229 941 348
rect 1081 364 1181 472
rect 1525 409 1625 515
rect 1801 482 1901 515
rect 1801 436 1814 482
rect 1860 449 1901 482
rect 2197 449 2297 515
rect 1860 436 2297 449
rect 1801 409 2297 436
rect 2421 426 2521 515
rect 1525 369 1753 409
rect 1081 351 1477 364
rect 1081 305 1418 351
rect 1464 305 1477 351
rect 1705 361 1753 369
rect 1705 348 2082 361
rect 1705 321 2023 348
rect 1081 292 1477 305
rect 1537 308 1657 321
rect 1081 232 1201 292
rect 1537 262 1598 308
rect 1644 262 1657 308
rect 1537 229 1657 262
rect 1781 302 2023 321
rect 2069 302 2082 348
rect 1781 289 2082 302
rect 1781 229 1901 289
rect 2177 229 2297 409
rect 2401 414 2521 426
rect 2401 368 2435 414
rect 2481 368 2521 414
rect 2401 229 2521 368
rect 2625 407 2725 515
rect 2829 471 2929 515
rect 3073 431 3173 515
rect 3073 412 3193 431
rect 2625 394 3017 407
rect 2625 348 2958 394
rect 3004 348 3017 394
rect 2849 335 3017 348
rect 3073 366 3106 412
rect 3152 366 3193 412
rect 2625 229 2745 288
rect 2849 229 2969 335
rect 3073 229 3193 366
rect 3297 355 3397 515
rect 3297 229 3417 355
rect 124 112 244 156
rect 348 112 468 156
rect 592 64 712 156
rect 821 112 941 156
rect 1081 112 1201 156
rect 1537 112 1657 156
rect 1781 112 1901 156
rect 2177 112 2297 156
rect 2401 112 2521 156
rect 2625 64 2745 156
rect 2849 112 2969 156
rect 3073 112 3193 156
rect 3297 64 3417 156
rect 592 24 3417 64
<< polycontact >>
rect 437 436 483 482
rect 141 348 187 394
rect 865 348 911 394
rect 653 262 699 308
rect 1814 436 1860 482
rect 1418 305 1464 351
rect 1598 262 1644 308
rect 2023 302 2069 348
rect 2435 368 2481 414
rect 2958 348 3004 394
rect 3106 366 3152 412
<< metal1 >>
rect 0 724 3584 844
rect 49 594 95 724
rect 527 620 906 666
rect 252 594 299 605
rect 527 594 595 620
rect 49 537 95 548
rect 141 394 202 590
rect 187 348 202 394
rect 49 215 95 226
rect 141 194 202 348
rect 252 548 253 594
rect 252 215 299 548
rect 345 548 538 594
rect 584 548 595 594
rect 345 314 391 548
rect 745 528 757 574
rect 803 528 814 574
rect 437 482 483 493
rect 437 424 483 436
rect 437 360 699 424
rect 345 268 458 314
rect 408 215 458 268
rect 640 308 699 360
rect 640 262 653 308
rect 640 248 699 262
rect 745 215 814 528
rect 860 523 906 620
rect 969 615 1037 724
rect 969 569 980 615
rect 1026 569 1037 615
rect 1104 631 1372 678
rect 1104 523 1150 631
rect 1326 601 1372 631
rect 1930 632 2271 678
rect 1326 590 1454 601
rect 1930 590 1976 632
rect 860 476 1150 523
rect 1198 525 1210 571
rect 1256 525 1276 571
rect 860 394 1110 430
rect 860 348 865 394
rect 911 360 1110 394
rect 911 348 917 360
rect 860 275 917 348
rect 1198 314 1276 525
rect 252 169 273 215
rect 319 169 330 215
rect 408 169 497 215
rect 543 169 554 215
rect 745 169 746 215
rect 792 169 814 215
rect 49 60 95 169
rect 745 156 814 169
rect 970 215 1016 232
rect 970 60 1016 169
rect 1130 215 1276 314
rect 1130 169 1230 215
rect 1130 120 1276 169
rect 1326 544 1408 590
rect 1326 533 1454 544
rect 1500 544 1694 590
rect 1740 544 1751 590
rect 1326 226 1372 533
rect 1500 364 1546 544
rect 1814 482 1860 493
rect 1814 430 1860 436
rect 1418 351 1546 364
rect 1464 305 1546 351
rect 1418 292 1546 305
rect 1326 215 1454 226
rect 1326 169 1405 215
rect 1451 169 1454 215
rect 1326 158 1454 169
rect 1500 152 1546 292
rect 1592 354 1860 430
rect 1592 308 1660 354
rect 1592 262 1598 308
rect 1644 262 1660 308
rect 1592 233 1660 262
rect 1706 215 1752 229
rect 1706 152 1752 169
rect 1930 215 1976 544
rect 1930 156 1976 169
rect 2022 574 2168 585
rect 2022 528 2122 574
rect 2022 515 2168 528
rect 2225 523 2271 632
rect 2334 615 2403 724
rect 2334 569 2346 615
rect 2392 569 2403 615
rect 2453 632 2820 678
rect 2453 523 2499 632
rect 2022 348 2070 515
rect 2225 476 2499 523
rect 2550 574 2596 585
rect 2118 414 2500 426
rect 2118 368 2435 414
rect 2481 368 2500 414
rect 2118 356 2500 368
rect 2022 302 2023 348
rect 2069 302 2070 348
rect 2022 229 2070 302
rect 2022 216 2168 229
rect 2022 170 2102 216
rect 2148 170 2168 216
rect 2022 159 2168 170
rect 2326 216 2372 229
rect 1500 106 1752 152
rect 2326 60 2372 170
rect 2550 216 2596 528
rect 2550 156 2596 170
rect 2754 574 2820 632
rect 3191 609 3259 724
rect 2800 528 2820 574
rect 2754 216 2820 528
rect 2754 170 2774 216
rect 2866 563 2981 609
rect 3027 563 3038 609
rect 3191 563 3202 609
rect 3248 563 3259 609
rect 3425 609 3492 628
rect 3425 563 3426 609
rect 3472 563 3492 609
rect 2866 216 2912 563
rect 3425 517 3492 563
rect 2958 471 3492 517
rect 2958 394 3004 471
rect 3050 412 3388 424
rect 3050 366 3106 412
rect 3152 366 3388 412
rect 3050 350 3388 366
rect 2958 337 3004 348
rect 3222 216 3268 229
rect 2866 170 2998 216
rect 3044 170 3055 216
rect 2754 156 2820 170
rect 3222 60 3268 170
rect 3446 216 3492 471
rect 3446 156 3492 170
rect 0 -60 3584 60
<< labels >>
flabel metal1 s 3050 350 3388 424 0 FreeSans 400 0 0 0 I0
port 1 nsew default input
flabel metal1 s 970 229 1016 232 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 0 724 3584 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 141 194 202 590 0 FreeSans 400 0 0 0 I2
port 3 nsew default input
flabel metal1 s 2118 356 2500 426 0 FreeSans 400 0 0 0 I1
port 2 nsew default input
flabel metal1 s 437 424 483 493 0 FreeSans 400 0 0 0 S0
port 5 nsew default input
flabel metal1 s 860 360 1110 430 0 FreeSans 400 0 0 0 I3
port 4 nsew default input
flabel metal1 s 1814 430 1860 493 0 FreeSans 400 0 0 0 S1
port 6 nsew default input
flabel metal1 s 1198 314 1276 571 0 FreeSans 400 0 0 0 Z
port 7 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 860 275 917 360 1 I3
port 4 nsew default input
rlabel metal1 s 437 360 699 424 1 S0
port 5 nsew default input
rlabel metal1 s 640 248 699 360 1 S0
port 5 nsew default input
rlabel metal1 s 1592 354 1860 430 1 S1
port 6 nsew default input
rlabel metal1 s 1592 233 1660 354 1 S1
port 6 nsew default input
rlabel metal1 s 1130 120 1276 314 1 Z
port 7 nsew default output
rlabel metal1 s 3191 569 3259 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2334 569 2403 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 969 569 1037 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 569 95 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3191 563 3259 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 563 95 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 537 95 563 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3222 226 3268 229 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 2326 226 2372 229 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 970 226 1016 229 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3222 60 3268 226 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 2326 60 2372 226 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 970 60 1016 226 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 226 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3584 60 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 784
string GDS_END 681862
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 673996
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
