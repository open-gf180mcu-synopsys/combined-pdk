magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 760 2045 830
rect 55 555 80 760
rect 55 518 105 520
rect 55 492 67 518
rect 93 492 105 518
rect 55 490 105 492
rect 385 630 410 760
rect 545 555 570 760
rect 850 555 875 760
rect 1130 630 1155 760
rect 340 453 390 455
rect 340 427 352 453
rect 378 427 390 453
rect 340 425 390 427
rect 595 388 645 390
rect 595 362 607 388
rect 633 362 645 388
rect 595 360 645 362
rect 55 70 80 190
rect 230 70 255 190
rect 1390 555 1415 760
rect 1550 680 1575 760
rect 1570 453 1620 455
rect 1570 427 1582 453
rect 1608 427 1620 453
rect 1570 425 1620 427
rect 455 70 480 190
rect 545 70 570 190
rect 850 70 875 150
rect 1130 70 1155 190
rect 1795 455 1820 725
rect 1880 555 1905 760
rect 1965 525 1990 725
rect 1965 518 2015 525
rect 1965 492 1977 518
rect 2003 492 2015 518
rect 1965 490 2015 492
rect 1965 485 2010 490
rect 1795 453 1940 455
rect 1795 427 1902 453
rect 1928 427 1940 453
rect 1795 425 1940 427
rect 1365 323 1415 325
rect 1365 297 1377 323
rect 1403 297 1415 323
rect 1365 295 1415 297
rect 1390 70 1415 190
rect 1480 70 1505 190
rect 1905 240 1930 425
rect 1795 215 1930 240
rect 1705 70 1730 190
rect 1795 105 1820 215
rect 1880 70 1905 190
rect 1965 105 1990 485
rect 0 0 2045 70
<< via1 >>
rect 67 492 93 518
rect 352 427 378 453
rect 607 362 633 388
rect 1582 427 1608 453
rect 1977 492 2003 518
rect 1902 427 1928 453
rect 1377 297 1403 323
<< obsm1 >>
rect 140 260 165 725
rect 215 285 240 725
rect 300 605 325 725
rect 470 605 495 725
rect 300 580 495 605
rect 710 530 735 725
rect 990 630 1015 725
rect 900 605 1015 630
rect 545 505 735 530
rect 545 390 570 505
rect 810 490 860 520
rect 665 425 780 455
rect 265 360 315 390
rect 440 360 570 390
rect 215 260 340 285
rect 450 260 475 265
rect 545 260 570 360
rect 740 260 770 425
rect 820 260 850 490
rect 900 380 925 605
rect 1075 490 1125 520
rect 1215 510 1240 725
rect 1305 565 1330 725
rect 895 355 925 380
rect 955 425 1060 455
rect 130 230 180 260
rect 315 230 490 260
rect 545 235 645 260
rect 140 225 170 230
rect 140 105 165 225
rect 315 105 340 230
rect 450 225 475 230
rect 605 190 645 235
rect 730 230 780 260
rect 810 230 860 260
rect 895 195 920 355
rect 955 255 985 425
rect 1085 390 1115 490
rect 1215 485 1270 510
rect 1170 425 1220 455
rect 1245 390 1270 485
rect 1300 455 1330 565
rect 1465 655 1490 725
rect 1635 655 1660 725
rect 1465 630 1660 655
rect 1480 520 1510 530
rect 1720 520 1745 725
rect 1480 490 1760 520
rect 1480 480 1510 490
rect 1295 425 1340 455
rect 1080 360 1130 390
rect 1215 365 1270 390
rect 1010 295 1060 325
rect 1215 285 1245 365
rect 945 225 995 255
rect 605 165 735 190
rect 895 170 1030 195
rect 710 105 735 165
rect 990 165 1030 170
rect 990 105 1015 165
rect 1215 105 1240 285
rect 1300 180 1330 425
rect 1720 325 1745 490
rect 1620 295 1865 325
rect 1470 225 1520 255
rect 1305 105 1330 180
rect 1620 105 1645 295
rect 1670 225 1720 255
<< metal2 >>
rect 350 555 1610 585
rect 55 518 105 525
rect 55 492 67 518
rect 93 492 105 518
rect 55 485 105 492
rect 350 460 380 555
rect 1580 460 1610 555
rect 1970 520 2010 525
rect 1965 518 2015 520
rect 1965 492 1977 518
rect 2003 492 2015 518
rect 1965 490 2015 492
rect 1970 485 2010 490
rect 340 453 390 460
rect 340 427 352 453
rect 378 427 390 453
rect 340 420 390 427
rect 1570 453 1620 460
rect 1895 455 1935 460
rect 1570 427 1582 453
rect 1608 427 1620 453
rect 1570 420 1620 427
rect 1890 453 1940 455
rect 1890 427 1902 453
rect 1928 427 1940 453
rect 1890 425 1940 427
rect 1895 420 1935 425
rect 595 388 645 395
rect 595 362 607 388
rect 633 362 645 388
rect 595 355 645 362
rect 1365 323 1415 330
rect 1365 297 1377 323
rect 1403 297 1415 323
rect 1365 290 1415 297
<< obsm2 >>
rect 1080 520 1120 525
rect 1475 520 1515 525
rect 1075 490 1520 520
rect 1080 485 1120 490
rect 1475 485 1515 490
rect 1710 485 1760 525
rect 730 455 775 460
rect 1010 455 1060 460
rect 1175 455 1215 460
rect 1295 455 1340 460
rect 730 425 1340 455
rect 730 420 775 425
rect 1010 420 1060 425
rect 1175 420 1215 425
rect 1295 420 1340 425
rect 265 355 315 395
rect 440 355 490 395
rect 1085 390 1125 395
rect 1080 360 1130 390
rect 1085 355 1125 360
rect 130 260 180 265
rect 275 260 305 355
rect 1015 325 1055 330
rect 1210 325 1250 330
rect 1010 295 1260 325
rect 1820 325 1860 330
rect 1015 290 1055 295
rect 1210 290 1250 295
rect 1785 295 1865 325
rect 1820 290 1860 295
rect 130 230 305 260
rect 130 225 180 230
rect 275 130 305 230
rect 440 260 490 265
rect 815 260 855 265
rect 440 230 860 260
rect 440 225 490 230
rect 815 225 855 230
rect 1470 220 1520 260
rect 1660 220 1720 260
rect 985 195 1025 200
rect 1470 195 1510 220
rect 980 165 1510 195
rect 985 160 1025 165
rect 1660 130 1690 220
rect 275 100 1690 130
<< labels >>
rlabel metal1 s 55 555 80 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 385 630 410 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 545 555 570 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 850 555 875 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1130 630 1155 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1390 555 1415 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1550 680 1575 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1880 555 1905 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 760 2045 830 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 55 0 80 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 230 0 255 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 455 0 480 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 545 0 570 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 850 0 875 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1130 0 1155 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1390 0 1415 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1480 0 1505 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1705 0 1730 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1880 0 1905 190 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2045 70 6 VSS
port 8 nsew ground bidirectional abutment
rlabel via1 s 1377 297 1403 323 6 CLK
port 4 nsew clock input
rlabel metal2 s 1365 290 1415 330 6 CLK
port 4 nsew clock input
rlabel metal1 s 1365 295 1415 325 6 CLK
port 4 nsew clock input
rlabel via1 s 607 362 633 388 6 D
port 1 nsew signal input
rlabel metal2 s 595 355 645 395 6 D
port 1 nsew signal input
rlabel metal1 s 595 360 645 390 6 D
port 1 nsew signal input
rlabel via1 s 1977 492 2003 518 6 Q
port 2 nsew signal output
rlabel metal2 s 1970 485 2010 525 6 Q
port 2 nsew signal output
rlabel metal2 s 1965 490 2015 520 6 Q
port 2 nsew signal output
rlabel metal1 s 1965 105 1990 725 6 Q
port 2 nsew signal output
rlabel metal1 s 1965 485 2010 525 6 Q
port 2 nsew signal output
rlabel metal1 s 1965 490 2015 525 6 Q
port 2 nsew signal output
rlabel via1 s 1902 427 1928 453 6 QN
port 3 nsew signal output
rlabel metal2 s 1895 420 1935 460 6 QN
port 3 nsew signal output
rlabel metal2 s 1890 425 1940 455 6 QN
port 3 nsew signal output
rlabel metal1 s 1795 105 1820 240 6 QN
port 3 nsew signal output
rlabel metal1 s 1795 425 1820 725 6 QN
port 3 nsew signal output
rlabel metal1 s 1795 215 1930 240 6 QN
port 3 nsew signal output
rlabel metal1 s 1905 215 1930 455 6 QN
port 3 nsew signal output
rlabel metal1 s 1795 425 1940 455 6 QN
port 3 nsew signal output
rlabel via1 s 67 492 93 518 6 RN
port 5 nsew signal input
rlabel metal2 s 55 485 105 525 6 RN
port 5 nsew signal input
rlabel metal1 s 55 490 105 520 6 RN
port 5 nsew signal input
rlabel via1 s 1582 427 1608 453 6 SN
port 6 nsew signal output
rlabel via1 s 352 427 378 453 6 SN
port 6 nsew signal output
rlabel metal2 s 350 420 380 585 6 SN
port 6 nsew signal output
rlabel metal2 s 340 420 390 460 6 SN
port 6 nsew signal output
rlabel metal2 s 1580 420 1610 585 6 SN
port 6 nsew signal output
rlabel metal2 s 350 555 1610 585 6 SN
port 6 nsew signal output
rlabel metal2 s 1570 420 1620 460 6 SN
port 6 nsew signal output
rlabel metal1 s 340 425 390 455 6 SN
port 6 nsew signal output
rlabel metal1 s 1570 425 1620 455 6 SN
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2045 830
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 375160
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 344958
<< end >>
