magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< isosubstrate >>
rect 2390 -6738 8471 -6737
rect 5759 -7815 8471 -6738
<< nwell >>
rect -83 53 8471 3035
rect 5925 -7651 7121 -6737
<< mvnmos >>
rect 7818 -7404 8118 -7264
<< mvpmos >>
rect 6278 -7404 6878 -7264
<< mvndiff >>
rect 7818 -7189 8118 -7176
rect 7818 -7235 7831 -7189
rect 7877 -7235 7945 -7189
rect 7991 -7235 8059 -7189
rect 8105 -7235 8118 -7189
rect 7818 -7264 8118 -7235
rect 7818 -7433 8118 -7404
rect 7818 -7479 7831 -7433
rect 7877 -7479 7945 -7433
rect 7991 -7479 8059 -7433
rect 8105 -7479 8118 -7433
rect 7818 -7492 8118 -7479
<< mvpdiff >>
rect 6278 -7189 6878 -7176
rect 6278 -7235 6291 -7189
rect 6337 -7235 6396 -7189
rect 6442 -7235 6501 -7189
rect 6547 -7235 6607 -7189
rect 6653 -7235 6713 -7189
rect 6759 -7235 6819 -7189
rect 6865 -7235 6878 -7189
rect 6278 -7264 6878 -7235
rect 6278 -7433 6878 -7404
rect 6278 -7479 6291 -7433
rect 6337 -7479 6396 -7433
rect 6442 -7479 6501 -7433
rect 6547 -7479 6607 -7433
rect 6653 -7479 6713 -7433
rect 6759 -7479 6819 -7433
rect 6865 -7479 6878 -7433
rect 6278 -7492 6878 -7479
<< mvndiffc >>
rect 7831 -7235 7877 -7189
rect 7945 -7235 7991 -7189
rect 8059 -7235 8105 -7189
rect 7831 -7479 7877 -7433
rect 7945 -7479 7991 -7433
rect 8059 -7479 8105 -7433
<< mvpdiffc >>
rect 6291 -7235 6337 -7189
rect 6396 -7235 6442 -7189
rect 6501 -7235 6547 -7189
rect 6607 -7235 6653 -7189
rect 6713 -7235 6759 -7189
rect 6819 -7235 6865 -7189
rect 6291 -7479 6337 -7433
rect 6396 -7479 6442 -7433
rect 6501 -7479 6547 -7433
rect 6607 -7479 6653 -7433
rect 6713 -7479 6759 -7433
rect 6819 -7479 6865 -7433
<< psubdiff >>
rect 7358 -6970 8388 -6948
rect 7358 -7016 7380 -6970
rect 8366 -7016 8388 -6970
rect 7358 -7038 8388 -7016
rect 8298 -7124 8388 -7038
rect 8298 -7546 8320 -7124
rect 8366 -7546 8388 -7124
rect 8298 -7632 8388 -7546
rect 7358 -7654 8388 -7632
rect 7358 -7700 7380 -7654
rect 8366 -7700 8388 -7654
rect 7358 -7722 8388 -7700
<< nsubdiff >>
rect 0 2930 8388 2952
rect 0 158 22 2930
rect 68 2884 176 2930
rect 8212 2884 8320 2930
rect 68 2862 8320 2884
rect 68 226 90 2862
rect 8298 2696 8320 2862
rect 8366 2696 8388 2930
rect 8298 2272 8388 2696
rect 8298 226 8320 2272
rect 68 204 8320 226
rect 68 158 176 204
rect 8212 158 8320 204
rect 8366 158 8388 2272
rect 0 136 8388 158
rect 6008 -6970 7038 -6948
rect 6008 -7016 6030 -6970
rect 7016 -7016 7038 -6970
rect 6008 -7038 7038 -7016
rect 6008 -7124 6098 -7038
rect 6008 -7546 6030 -7124
rect 6076 -7546 6098 -7124
rect 6008 -7568 6098 -7546
<< psubdiffcont >>
rect 7380 -7016 8366 -6970
rect 8320 -7546 8366 -7124
rect 7380 -7700 8366 -7654
<< nsubdiffcont >>
rect 22 158 68 2930
rect 176 2884 8212 2930
rect 8320 2696 8366 2930
rect 176 158 8212 204
rect 8320 158 8366 2272
rect 6030 -7016 7016 -6970
rect 6030 -7546 6076 -7124
<< polysilicon >>
rect 404 2547 506 2604
rect 404 2501 417 2547
rect 463 2501 506 2547
rect 404 2444 506 2501
rect 7646 2547 7748 2604
rect 7646 2501 7689 2547
rect 7735 2501 7748 2547
rect 7646 2444 7748 2501
rect 404 2267 506 2324
rect 404 2221 417 2267
rect 463 2221 506 2267
rect 404 2164 506 2221
rect 7646 2267 7748 2324
rect 7646 2221 7689 2267
rect 7735 2221 7748 2267
rect 7646 2164 7748 2221
rect 404 1987 506 2044
rect 404 1941 417 1987
rect 463 1941 506 1987
rect 404 1884 506 1941
rect 7646 1987 7748 2044
rect 7646 1941 7689 1987
rect 7735 1941 7748 1987
rect 7646 1884 7748 1941
rect 404 1707 506 1764
rect 404 1661 417 1707
rect 463 1661 506 1707
rect 404 1604 506 1661
rect 7646 1707 7748 1764
rect 7646 1661 7689 1707
rect 7735 1661 7748 1707
rect 7646 1604 7748 1661
rect 404 1427 506 1484
rect 404 1381 417 1427
rect 463 1381 506 1427
rect 404 1324 506 1381
rect 7646 1427 7748 1484
rect 7646 1381 7689 1427
rect 7735 1381 7748 1427
rect 7646 1324 7748 1381
rect 404 1147 506 1204
rect 404 1101 417 1147
rect 463 1101 506 1147
rect 404 1044 506 1101
rect 7646 1147 7748 1204
rect 7646 1101 7689 1147
rect 7735 1101 7748 1147
rect 7646 1044 7748 1101
rect 404 867 506 924
rect 404 821 417 867
rect 463 821 506 867
rect 404 764 506 821
rect 7646 867 7748 924
rect 7646 821 7689 867
rect 7735 821 7748 867
rect 7646 764 7748 821
rect 404 587 506 644
rect 404 541 417 587
rect 463 541 506 587
rect 404 484 506 541
rect 5106 587 5208 644
rect 5106 541 5149 587
rect 5195 541 5208 587
rect 5106 484 5208 541
rect 6234 -7404 6278 -7264
rect 6878 -7311 7092 -7264
rect 6878 -7357 6933 -7311
rect 7073 -7357 7092 -7311
rect 6878 -7404 7092 -7357
rect 7477 -7311 7818 -7264
rect 7477 -7357 7496 -7311
rect 7636 -7357 7818 -7311
rect 7477 -7404 7818 -7357
rect 8118 -7404 8162 -7264
<< polycontact >>
rect 417 2501 463 2547
rect 7689 2501 7735 2547
rect 417 2221 463 2267
rect 7689 2221 7735 2267
rect 417 1941 463 1987
rect 7689 1941 7735 1987
rect 417 1661 463 1707
rect 7689 1661 7735 1707
rect 417 1381 463 1427
rect 7689 1381 7735 1427
rect 417 1101 463 1147
rect 7689 1101 7735 1147
rect 417 821 463 867
rect 7689 821 7735 867
rect 417 541 463 587
rect 5149 541 5195 587
rect 6933 -7357 7073 -7311
rect 7496 -7357 7636 -7311
<< ppolyres >>
rect 506 2444 7646 2604
rect 506 2164 7646 2324
rect 506 1884 7646 2044
rect 506 1604 7646 1764
rect 506 1324 7646 1484
rect 506 1044 7646 1204
rect 506 764 7646 924
rect 506 484 5106 644
<< metal1 >>
rect 11 2930 8377 2941
rect 11 158 22 2930
rect 68 2884 176 2930
rect 8212 2884 8320 2930
rect 68 2873 8320 2884
rect 68 215 79 2873
rect 8309 2696 8320 2873
rect 8366 2696 8377 2930
rect 8309 2669 8377 2696
rect 406 2547 474 2602
rect 406 2501 417 2547
rect 463 2501 474 2547
rect 406 2267 474 2501
rect 7678 2547 8992 2602
rect 7678 2501 7689 2547
rect 7735 2501 8992 2547
rect 7678 2446 8992 2501
rect 406 2221 417 2267
rect 463 2221 474 2267
rect 406 2166 474 2221
rect 7678 2267 7746 2322
rect 7678 2221 7689 2267
rect 7735 2221 7746 2267
rect 406 1987 474 2042
rect 406 1941 417 1987
rect 463 1941 474 1987
rect 406 1707 474 1941
rect 7678 1987 7746 2221
rect 7678 1941 7689 1987
rect 7735 1941 7746 1987
rect 7678 1886 7746 1941
rect 8309 2272 8377 2338
rect 406 1661 417 1707
rect 463 1661 474 1707
rect 406 1606 474 1661
rect 7678 1707 7746 1762
rect 7678 1661 7689 1707
rect 7735 1661 7746 1707
rect 406 1427 474 1482
rect 406 1381 417 1427
rect 463 1381 474 1427
rect 406 1147 474 1381
rect 7678 1427 7746 1661
rect 7678 1381 7689 1427
rect 7735 1381 7746 1427
rect 7678 1326 7746 1381
rect 406 1101 417 1147
rect 463 1101 474 1147
rect 406 1046 474 1101
rect 7678 1147 7746 1202
rect 7678 1101 7689 1147
rect 7735 1101 7746 1147
rect 406 867 474 922
rect 406 821 417 867
rect 463 821 474 867
rect 406 587 474 821
rect 7678 867 7746 1101
rect 7678 821 7689 867
rect 7735 821 7746 867
rect 7678 766 7746 821
rect 406 541 417 587
rect 463 541 474 587
rect 406 486 474 541
rect 5138 587 5206 642
rect 5138 541 5149 587
rect 5195 541 5206 587
rect 5138 486 5206 541
rect 8309 215 8320 2272
rect 68 204 8320 215
rect 68 158 176 204
rect 8212 158 8320 204
rect 8366 158 8377 2272
rect 11 147 8377 158
rect 6019 -6970 7027 -6959
rect 6019 -7016 6030 -6970
rect 7016 -7016 7027 -6970
rect 6019 -7027 7027 -7016
rect 7369 -6970 8377 -6959
rect 7369 -7016 7380 -6970
rect 8366 -7016 8377 -6970
rect 7369 -7027 8377 -7016
rect 6019 -7124 6087 -7027
rect 6019 -7546 6030 -7124
rect 6076 -7174 6087 -7124
rect 8309 -7124 8377 -7027
rect 8309 -7174 8320 -7124
rect 6076 -7189 6878 -7174
rect 6076 -7235 6291 -7189
rect 6337 -7235 6396 -7189
rect 6442 -7235 6501 -7189
rect 6547 -7235 6607 -7189
rect 6653 -7235 6713 -7189
rect 6759 -7235 6819 -7189
rect 6865 -7235 6878 -7189
rect 6076 -7250 6878 -7235
rect 7818 -7189 8320 -7174
rect 7818 -7235 7831 -7189
rect 7877 -7235 7945 -7189
rect 7991 -7235 8059 -7189
rect 8105 -7235 8320 -7189
rect 7818 -7250 8320 -7235
rect 6076 -7546 6087 -7250
rect 6922 -7311 7084 -7300
rect 6922 -7357 6933 -7311
rect 7073 -7357 7084 -7311
rect 6922 -7368 7084 -7357
rect 7485 -7311 7647 -7300
rect 7485 -7357 7496 -7311
rect 7636 -7357 7647 -7311
rect 7485 -7368 7647 -7357
rect 6278 -7433 8118 -7418
rect 6278 -7479 6291 -7433
rect 6337 -7479 6396 -7433
rect 6442 -7479 6501 -7433
rect 6547 -7479 6607 -7433
rect 6653 -7479 6713 -7433
rect 6759 -7479 6819 -7433
rect 6865 -7479 7831 -7433
rect 7877 -7479 7945 -7433
rect 7991 -7452 8059 -7433
rect 8105 -7452 8118 -7433
rect 6278 -7494 7950 -7479
rect 7938 -7504 7950 -7494
rect 8106 -7504 8118 -7452
rect 7938 -7516 8118 -7504
rect 6019 -7557 6087 -7546
rect 8309 -7546 8320 -7250
rect 8366 -7546 8377 -7124
rect 8836 -7440 8992 2446
rect 8812 -7452 8992 -7440
rect 8812 -7504 8824 -7452
rect 8980 -7504 8992 -7452
rect 8812 -7516 8992 -7504
rect 8309 -7643 8377 -7546
rect 7369 -7654 8377 -7643
rect 7369 -7700 7380 -7654
rect 8366 -7700 8377 -7654
rect 7369 -7711 8377 -7700
<< via1 >>
rect 7950 -7479 7991 -7452
rect 7991 -7479 8059 -7452
rect 8059 -7479 8105 -7452
rect 8105 -7479 8106 -7452
rect 7950 -7504 8106 -7479
rect 8824 -7504 8980 -7452
<< metal2 >>
rect 7938 -7452 8992 -7440
rect 7938 -7504 7950 -7452
rect 8106 -7504 8824 -7452
rect 8980 -7504 8992 -7452
rect 7938 -7516 8992 -7504
use M1_NWELL_CDNS_40661956134335  M1_NWELL_CDNS_40661956134335_0
timestamp 1750858719
transform 1 0 45 0 -1 1544
box 0 0 1 1
use M1_NWELL_CDNS_40661956134377  M1_NWELL_CDNS_40661956134377_0
timestamp 1750858719
transform 0 -1 6053 -1 0 -7335
box 0 0 1 1
use M1_NWELL_CDNS_40661956134418  M1_NWELL_CDNS_40661956134418_0
timestamp 1750858719
transform 0 -1 6523 -1 0 -6993
box 0 0 1 1
use M1_NWELL_CDNS_40661956134419  M1_NWELL_CDNS_40661956134419_0
timestamp 1750858719
transform 1 0 4194 0 -1 181
box 0 0 1 1
use M1_NWELL_CDNS_40661956134419  M1_NWELL_CDNS_40661956134419_1
timestamp 1750858719
transform 1 0 4194 0 -1 2907
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_0
timestamp 1750858719
transform 0 -1 7566 1 0 -7334
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_1
timestamp 1750858719
transform 0 -1 7003 1 0 -7334
box 0 0 1 1
use M1_PSUB_CDNS_40661956134330  M1_PSUB_CDNS_40661956134330_0
timestamp 1750858719
transform 0 1 7873 -1 0 -6993
box 0 0 1 1
use M1_PSUB_CDNS_40661956134330  M1_PSUB_CDNS_40661956134330_1
timestamp 1750858719
transform 0 1 7873 -1 0 -7677
box 0 0 1 1
use M1_PSUB_CDNS_40661956134341  M1_PSUB_CDNS_40661956134341_0
timestamp 1750858719
transform 0 1 8343 -1 0 -7335
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_0
timestamp 1750858719
transform 1 0 8028 0 1 -7478
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_1
timestamp 1750858719
transform 1 0 8902 0 1 -7478
box 0 0 1 1
use nmos_6p0_CDNS_4066195613430  nmos_6p0_CDNS_4066195613430_0
timestamp 1750858719
transform 0 -1 8118 -1 0 -7264
box 0 0 1 1
use pmos_6p0_CDNS_4066195613412  pmos_6p0_CDNS_4066195613412_0
timestamp 1750858719
transform 0 -1 6878 -1 0 -7264
box 0 0 1 1
use ppolyf_u_CDNS_4066195613432  ppolyf_u_CDNS_4066195613432_0
timestamp 1750858719
transform -1 0 5208 0 1 484
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_0
timestamp 1750858719
transform -1 0 7748 0 1 1604
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_1
timestamp 1750858719
transform -1 0 7748 0 1 1044
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_2
timestamp 1750858719
transform 1 0 404 0 1 2444
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_3
timestamp 1750858719
transform 1 0 404 0 1 2164
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_4
timestamp 1750858719
transform 1 0 404 0 1 1884
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_5
timestamp 1750858719
transform 1 0 404 0 1 1324
box 0 0 1 1
use ppolyf_u_CDNS_4066195613433  ppolyf_u_CDNS_4066195613433_6
timestamp 1750858719
transform 1 0 404 0 1 764
box 0 0 1 1
<< labels >>
rlabel metal1 s 5175 575 5175 575 4 A
port 1 nsew
rlabel metal1 s 6048 -7005 6048 -7005 4 DVDD
port 2 nsew
rlabel metal1 s 8343 -7192 8343 -7192 4 DVSS
port 3 nsew
rlabel metal1 s 7110 -7333 7110 -7333 4 PU_B
port 4 nsew
rlabel metal1 s 7561 -7333 7561 -7333 4 PD
port 5 nsew
<< properties >>
string GDS_END 989476
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 983576
string path 224.800 -186.950 198.450 -186.950 
<< end >>
