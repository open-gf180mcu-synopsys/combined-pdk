magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 780 1660
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
rect 500 210 560 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 530 1110 590 1450
<< ndiff >>
rect 120 318 220 380
rect 120 272 142 318
rect 188 272 220 318
rect 120 210 220 272
rect 280 210 330 380
rect 390 318 500 380
rect 390 272 422 318
rect 468 272 500 318
rect 390 210 500 272
rect 560 318 660 380
rect 560 272 592 318
rect 638 272 660 318
rect 560 210 660 272
<< pdiff >>
rect 90 1425 190 1450
rect 90 1285 112 1425
rect 158 1285 190 1425
rect 90 1110 190 1285
rect 250 1425 360 1450
rect 250 1285 282 1425
rect 328 1285 360 1425
rect 250 1110 360 1285
rect 420 1425 530 1450
rect 420 1285 452 1425
rect 498 1285 530 1425
rect 420 1110 530 1285
rect 590 1397 690 1450
rect 590 1163 622 1397
rect 668 1163 690 1397
rect 590 1110 690 1163
<< ndiffc >>
rect 142 272 188 318
rect 422 272 468 318
rect 592 272 638 318
<< pdiffc >>
rect 112 1285 158 1425
rect 282 1285 328 1425
rect 452 1285 498 1425
rect 622 1163 668 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 530 1450 590 1500
rect 190 800 250 1110
rect 360 930 420 1110
rect 300 903 420 930
rect 300 857 347 903
rect 393 857 420 903
rect 300 830 420 857
rect 110 773 250 800
rect 110 727 147 773
rect 193 727 250 773
rect 110 700 250 727
rect 190 470 250 700
rect 360 470 420 830
rect 530 800 590 1110
rect 470 773 590 800
rect 470 727 497 773
rect 543 727 590 773
rect 470 700 590 727
rect 530 650 590 700
rect 190 430 280 470
rect 220 380 280 430
rect 330 430 420 470
rect 500 610 590 650
rect 330 380 390 430
rect 500 380 560 610
rect 220 160 280 210
rect 330 160 390 210
rect 500 160 560 210
<< polycontact >>
rect 347 857 393 903
rect 147 727 193 773
rect 497 727 543 773
<< metal1 >>
rect 0 1588 780 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 780 1588
rect 0 1520 780 1542
rect 110 1425 160 1450
rect 110 1285 112 1425
rect 158 1285 160 1425
rect 110 1210 160 1285
rect 280 1425 330 1520
rect 280 1285 282 1425
rect 328 1285 330 1425
rect 280 1260 330 1285
rect 450 1425 500 1450
rect 450 1285 452 1425
rect 498 1285 500 1425
rect 450 1210 500 1285
rect 110 1160 500 1210
rect 620 1397 670 1450
rect 620 1163 622 1397
rect 668 1163 670 1397
rect 620 1040 670 1163
rect 600 1036 700 1040
rect 600 984 624 1036
rect 676 984 700 1036
rect 600 980 700 984
rect 320 906 420 910
rect 320 854 344 906
rect 396 854 420 906
rect 320 850 420 854
rect 120 776 220 780
rect 120 724 144 776
rect 196 724 220 776
rect 120 720 220 724
rect 470 776 570 780
rect 470 724 494 776
rect 546 724 570 776
rect 470 720 570 724
rect 620 580 670 980
rect 420 530 670 580
rect 140 318 190 380
rect 140 272 142 318
rect 188 272 190 318
rect 140 140 190 272
rect 420 318 470 530
rect 420 272 422 318
rect 468 272 470 318
rect 420 210 470 272
rect 590 318 640 380
rect 590 272 592 318
rect 638 272 640 318
rect 590 140 640 272
rect 0 118 780 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 780 118
rect 0 0 780 72
<< via1 >>
rect 624 984 676 1036
rect 344 903 396 906
rect 344 857 347 903
rect 347 857 393 903
rect 393 857 396 903
rect 344 854 396 857
rect 144 773 196 776
rect 144 727 147 773
rect 147 727 193 773
rect 193 727 196 773
rect 144 724 196 727
rect 494 773 546 776
rect 494 727 497 773
rect 497 727 543 773
rect 543 727 546 773
rect 494 724 546 727
<< metal2 >>
rect 600 1036 700 1050
rect 600 984 624 1036
rect 676 984 700 1036
rect 600 970 700 984
rect 320 906 420 920
rect 320 854 344 906
rect 396 854 420 906
rect 320 840 420 854
rect 120 776 220 790
rect 120 724 144 776
rect 196 724 220 776
rect 120 710 220 724
rect 470 776 570 790
rect 470 724 494 776
rect 546 724 570 776
rect 470 710 570 724
<< labels >>
rlabel via1 s 144 724 196 776 4 A0
port 1 nsew signal input
rlabel via1 s 344 854 396 906 4 A1
port 2 nsew signal input
rlabel via1 s 494 724 546 776 4 B
port 3 nsew signal input
rlabel via1 s 624 984 676 1036 4 Y
port 4 nsew signal output
rlabel metal1 s 280 1260 330 1660 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 140 0 190 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 1520 780 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 590 0 640 380 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 780 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 120 710 220 790 1 A0
port 1 nsew signal input
rlabel metal1 s 120 720 220 780 1 A0
port 1 nsew signal input
rlabel metal2 s 320 840 420 920 1 A1
port 2 nsew signal input
rlabel metal1 s 320 850 420 910 1 A1
port 2 nsew signal input
rlabel metal2 s 470 710 570 790 1 B
port 3 nsew signal input
rlabel metal1 s 470 720 570 780 1 B
port 3 nsew signal input
rlabel metal2 s 600 970 700 1050 1 Y
port 4 nsew signal output
rlabel metal1 s 420 210 470 580 1 Y
port 4 nsew signal output
rlabel metal1 s 420 530 670 580 1 Y
port 4 nsew signal output
rlabel metal1 s 620 530 670 1450 1 Y
port 4 nsew signal output
rlabel metal1 s 600 980 700 1040 1 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 780 1660
string GDS_END 41348
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 35928
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
