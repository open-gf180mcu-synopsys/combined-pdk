magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 1040 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 470 210 530 380
rect 790 210 850 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 470 1110 530 1450
rect 790 1110 850 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 470 380
rect 530 318 630 380
rect 530 272 562 318
rect 608 272 630 318
rect 530 210 630 272
rect 690 318 790 380
rect 690 272 712 318
rect 758 272 790 318
rect 690 210 790 272
rect 850 318 950 380
rect 850 272 882 318
rect 928 272 950 318
rect 850 210 950 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1110 470 1450
rect 530 1397 630 1450
rect 530 1163 562 1397
rect 608 1163 630 1397
rect 530 1110 630 1163
rect 690 1397 790 1450
rect 690 1163 712 1397
rect 758 1163 790 1397
rect 690 1110 790 1163
rect 850 1397 950 1450
rect 850 1163 882 1397
rect 928 1163 950 1397
rect 850 1110 950 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 562 272 608 318
rect 712 272 758 318
rect 882 272 928 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 562 1163 608 1397
rect 712 1163 758 1397
rect 882 1163 928 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 470 1450 530 1500
rect 790 1450 850 1500
rect 190 930 250 1110
rect 190 903 310 930
rect 190 857 237 903
rect 283 857 310 903
rect 190 830 310 857
rect 190 380 250 830
rect 360 780 420 1110
rect 470 1050 530 1110
rect 470 1028 580 1050
rect 470 982 512 1028
rect 558 982 580 1028
rect 470 960 580 982
rect 300 743 420 780
rect 300 697 327 743
rect 373 697 420 743
rect 300 660 420 697
rect 360 380 420 660
rect 600 518 700 540
rect 600 510 622 518
rect 470 472 622 510
rect 668 510 700 518
rect 790 510 850 1110
rect 668 472 850 510
rect 470 450 850 472
rect 470 380 530 450
rect 790 380 850 450
rect 190 160 250 210
rect 360 160 420 210
rect 470 160 530 210
rect 790 160 850 210
<< polycontact >>
rect 237 857 283 903
rect 512 982 558 1028
rect 327 697 373 743
rect 622 472 668 518
<< metal1 >>
rect 0 1588 1040 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1040 1588
rect 0 1520 1040 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 750 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 560 1397 610 1450
rect 560 1163 562 1397
rect 608 1163 610 1397
rect 560 1160 610 1163
rect 390 1110 610 1160
rect 710 1397 760 1520
rect 710 1163 712 1397
rect 758 1163 760 1397
rect 710 1110 760 1163
rect 880 1397 930 1450
rect 880 1163 882 1397
rect 928 1163 930 1397
rect 390 920 440 1110
rect 880 1040 930 1163
rect 490 1036 590 1040
rect 490 1028 514 1036
rect 490 982 512 1028
rect 566 984 590 1036
rect 558 982 590 984
rect 490 980 590 982
rect 860 1036 960 1040
rect 860 984 884 1036
rect 936 984 960 1036
rect 860 980 960 984
rect 210 906 310 910
rect 210 854 234 906
rect 286 854 310 906
rect 390 870 560 920
rect 210 850 310 854
rect 510 780 560 870
rect 490 776 590 780
rect 110 743 400 750
rect 110 697 327 743
rect 373 697 400 743
rect 490 724 514 776
rect 566 724 590 776
rect 490 720 590 724
rect 110 690 400 697
rect 110 318 160 690
rect 510 620 560 720
rect 390 570 560 620
rect 390 380 440 570
rect 600 526 700 530
rect 600 518 624 526
rect 600 472 622 518
rect 676 474 700 526
rect 668 472 700 474
rect 600 470 700 472
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 390 330 610 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 560 318 610 330
rect 560 272 562 318
rect 608 272 610 318
rect 560 210 610 272
rect 710 318 760 380
rect 710 272 712 318
rect 758 272 760 318
rect 710 140 760 272
rect 880 318 930 980
rect 880 272 882 318
rect 928 272 930 318
rect 880 210 930 272
rect 0 118 1040 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1040 118
rect 0 0 1040 72
<< via1 >>
rect 514 1028 566 1036
rect 514 984 558 1028
rect 558 984 566 1028
rect 884 984 936 1036
rect 234 903 286 906
rect 234 857 237 903
rect 237 857 283 903
rect 283 857 286 903
rect 234 854 286 857
rect 514 724 566 776
rect 624 518 676 526
rect 624 474 668 518
rect 668 474 676 518
<< metal2 >>
rect 490 1040 590 1050
rect 860 1040 960 1050
rect 490 1036 960 1040
rect 490 984 514 1036
rect 566 984 884 1036
rect 936 984 960 1036
rect 490 980 960 984
rect 490 970 590 980
rect 860 970 960 980
rect 220 910 300 920
rect 210 906 310 910
rect 210 854 234 906
rect 286 854 310 906
rect 210 850 310 854
rect 220 840 300 850
rect 490 776 590 790
rect 490 724 514 776
rect 566 724 590 776
rect 490 710 590 724
rect 600 526 700 540
rect 600 474 624 526
rect 676 474 700 526
rect 600 460 700 474
<< labels >>
rlabel via1 s 234 854 286 906 4 A
port 1 nsew signal input
rlabel via1 s 514 724 566 776 4 Y
port 2 nsew signal output
rlabel via1 s 624 474 676 526 4 EN
port 3 nsew signal input
rlabel metal1 s 280 1110 330 1660 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 710 1110 760 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1520 1040 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 710 0 760 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1040 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 220 840 300 920 1 A
port 1 nsew signal input
rlabel metal2 s 210 850 310 910 1 A
port 1 nsew signal input
rlabel metal1 s 210 850 310 910 1 A
port 1 nsew signal input
rlabel metal2 s 600 460 700 540 1 EN
port 3 nsew signal input
rlabel metal1 s 600 470 700 530 1 EN
port 3 nsew signal input
rlabel metal2 s 490 710 590 790 1 Y
port 2 nsew signal output
rlabel metal1 s 390 330 440 620 1 Y
port 2 nsew signal output
rlabel metal1 s 390 870 440 1160 1 Y
port 2 nsew signal output
rlabel metal1 s 390 570 560 620 1 Y
port 2 nsew signal output
rlabel metal1 s 390 1110 610 1160 1 Y
port 2 nsew signal output
rlabel metal1 s 510 570 560 920 1 Y
port 2 nsew signal output
rlabel metal1 s 390 870 560 920 1 Y
port 2 nsew signal output
rlabel metal1 s 490 720 590 780 1 Y
port 2 nsew signal output
rlabel metal1 s 560 210 610 380 1 Y
port 2 nsew signal output
rlabel metal1 s 390 330 610 380 1 Y
port 2 nsew signal output
rlabel metal1 s 560 1110 610 1450 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1040 1660
string GDS_END 504516
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 497214
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
