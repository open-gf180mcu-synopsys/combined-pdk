magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 982 1094
<< pwell >>
rect -86 -86 982 453
<< metal1 >>
rect 0 918 896 1098
rect 49 710 95 918
rect 273 664 319 872
rect 477 710 523 918
rect 701 664 747 872
rect 273 618 747 664
rect 82 454 432 542
rect 478 390 561 618
rect 273 344 767 390
rect 49 90 95 298
rect 273 136 319 344
rect 497 90 543 298
rect 721 136 767 344
rect 0 -90 896 90
<< labels >>
rlabel metal1 s 82 454 432 542 6 I
port 1 nsew default input
rlabel metal1 s 721 136 767 344 6 ZN
port 2 nsew default output
rlabel metal1 s 273 136 319 344 6 ZN
port 2 nsew default output
rlabel metal1 s 273 344 767 390 6 ZN
port 2 nsew default output
rlabel metal1 s 478 390 561 618 6 ZN
port 2 nsew default output
rlabel metal1 s 273 618 747 664 6 ZN
port 2 nsew default output
rlabel metal1 s 701 664 747 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 664 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 477 710 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 896 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 982 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 982 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 896 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 877472
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 874154
<< end >>
