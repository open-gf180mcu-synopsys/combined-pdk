magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 2800 1670
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
rect 870 210 930 380
rect 1040 210 1100 380
rect 1210 210 1270 380
rect 1380 210 1440 380
rect 1550 210 1610 380
rect 1720 210 1780 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2550 210 2610 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 530 1110 590 1450
rect 700 1110 760 1450
rect 870 1110 930 1450
rect 1040 1110 1100 1450
rect 1210 1110 1270 1450
rect 1380 1110 1440 1450
rect 1550 1110 1610 1450
rect 1720 1110 1780 1450
rect 1890 1110 1950 1450
rect 2060 1110 2120 1450
rect 2230 1110 2290 1450
rect 2550 1110 2610 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 318 530 380
rect 420 272 452 318
rect 498 272 530 318
rect 420 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 210 870 380
rect 930 318 1040 380
rect 930 272 962 318
rect 1008 272 1040 318
rect 930 210 1040 272
rect 1100 313 1210 380
rect 1100 267 1132 313
rect 1178 267 1210 313
rect 1100 210 1210 267
rect 1270 283 1380 380
rect 1270 237 1302 283
rect 1348 237 1380 283
rect 1270 210 1380 237
rect 1440 313 1550 380
rect 1440 267 1472 313
rect 1518 267 1550 313
rect 1440 210 1550 267
rect 1610 318 1720 380
rect 1610 272 1642 318
rect 1688 272 1720 318
rect 1610 210 1720 272
rect 1780 210 1890 380
rect 1950 210 2060 380
rect 2120 318 2230 380
rect 2120 272 2152 318
rect 2198 272 2230 318
rect 2120 210 2230 272
rect 2290 318 2390 380
rect 2290 272 2322 318
rect 2368 272 2390 318
rect 2290 210 2390 272
rect 2450 318 2550 380
rect 2450 272 2472 318
rect 2518 272 2550 318
rect 2450 210 2550 272
rect 2610 318 2710 380
rect 2610 272 2642 318
rect 2688 272 2710 318
rect 2610 210 2710 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1397 530 1450
rect 420 1163 452 1397
rect 498 1163 530 1397
rect 420 1110 530 1163
rect 590 1397 700 1450
rect 590 1163 622 1397
rect 668 1163 700 1397
rect 590 1110 700 1163
rect 760 1110 870 1450
rect 930 1397 1040 1450
rect 930 1163 962 1397
rect 1008 1163 1040 1397
rect 930 1110 1040 1163
rect 1100 1397 1210 1450
rect 1100 1163 1132 1397
rect 1178 1163 1210 1397
rect 1100 1110 1210 1163
rect 1270 1397 1380 1450
rect 1270 1163 1302 1397
rect 1348 1163 1380 1397
rect 1270 1110 1380 1163
rect 1440 1397 1550 1450
rect 1440 1163 1472 1397
rect 1518 1163 1550 1397
rect 1440 1110 1550 1163
rect 1610 1397 1720 1450
rect 1610 1163 1642 1397
rect 1688 1163 1720 1397
rect 1610 1110 1720 1163
rect 1780 1110 1890 1450
rect 1950 1110 2060 1450
rect 2120 1397 2230 1450
rect 2120 1163 2152 1397
rect 2198 1163 2230 1397
rect 2120 1110 2230 1163
rect 2290 1397 2390 1450
rect 2290 1163 2322 1397
rect 2368 1163 2390 1397
rect 2290 1110 2390 1163
rect 2450 1397 2550 1450
rect 2450 1163 2472 1397
rect 2518 1163 2550 1397
rect 2450 1110 2550 1163
rect 2610 1397 2710 1450
rect 2610 1163 2642 1397
rect 2688 1163 2710 1397
rect 2610 1110 2710 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 962 272 1008 318
rect 1132 267 1178 313
rect 1302 237 1348 283
rect 1472 267 1518 313
rect 1642 272 1688 318
rect 2152 272 2198 318
rect 2322 272 2368 318
rect 2472 272 2518 318
rect 2642 272 2688 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 452 1163 498 1397
rect 622 1163 668 1397
rect 962 1163 1008 1397
rect 1132 1163 1178 1397
rect 1302 1163 1348 1397
rect 1472 1163 1518 1397
rect 1642 1163 1688 1397
rect 2152 1163 2198 1397
rect 2322 1163 2368 1397
rect 2472 1163 2518 1397
rect 2642 1163 2688 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1020 1588 1170 1610
rect 1020 1542 1072 1588
rect 1118 1542 1170 1588
rect 1020 1520 1170 1542
rect 1260 1588 1410 1610
rect 1260 1542 1312 1588
rect 1358 1542 1410 1588
rect 1260 1520 1410 1542
rect 1500 1588 1650 1610
rect 1500 1542 1552 1588
rect 1598 1542 1650 1588
rect 1500 1520 1650 1542
rect 1740 1588 1890 1610
rect 1740 1542 1792 1588
rect 1838 1542 1890 1588
rect 1740 1520 1890 1542
rect 1980 1588 2130 1610
rect 1980 1542 2032 1588
rect 2078 1542 2130 1588
rect 1980 1520 2130 1542
rect 2220 1588 2370 1610
rect 2220 1542 2272 1588
rect 2318 1542 2370 1588
rect 2220 1520 2370 1542
rect 2460 1588 2610 1610
rect 2460 1542 2512 1588
rect 2558 1542 2610 1588
rect 2460 1520 2610 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1072 1542 1118 1588
rect 1312 1542 1358 1588
rect 1552 1542 1598 1588
rect 1792 1542 1838 1588
rect 2032 1542 2078 1588
rect 2272 1542 2318 1588
rect 2512 1542 2558 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 530 1450 590 1500
rect 700 1450 760 1500
rect 870 1450 930 1500
rect 1040 1450 1100 1500
rect 1210 1450 1270 1500
rect 1380 1450 1440 1500
rect 1550 1450 1610 1500
rect 1720 1450 1780 1500
rect 1890 1450 1950 1500
rect 2060 1450 2120 1500
rect 2230 1450 2290 1500
rect 2550 1450 2610 1500
rect 190 800 250 1110
rect 360 930 420 1110
rect 300 903 420 930
rect 300 857 327 903
rect 373 857 420 903
rect 300 830 420 857
rect 120 773 250 800
rect 120 727 147 773
rect 193 727 250 773
rect 120 700 250 727
rect 190 380 250 700
rect 360 380 420 830
rect 530 670 590 1110
rect 470 643 590 670
rect 470 597 497 643
rect 543 597 590 643
rect 470 570 590 597
rect 530 380 590 570
rect 700 930 760 1110
rect 870 1090 930 1110
rect 1040 1090 1100 1110
rect 870 1040 1100 1090
rect 700 903 820 930
rect 700 857 747 903
rect 793 857 820 903
rect 700 830 820 857
rect 700 380 760 830
rect 870 800 930 1040
rect 1210 930 1270 1110
rect 1150 903 1270 930
rect 1150 857 1177 903
rect 1223 857 1270 903
rect 1150 830 1270 857
rect 870 773 1020 800
rect 870 727 947 773
rect 993 727 1020 773
rect 870 700 1020 727
rect 870 450 930 700
rect 870 400 1100 450
rect 870 380 930 400
rect 1040 380 1100 400
rect 1210 380 1270 830
rect 1380 540 1440 1110
rect 1550 670 1610 1110
rect 1490 643 1610 670
rect 1490 597 1517 643
rect 1563 597 1610 643
rect 1490 570 1610 597
rect 1330 513 1440 540
rect 1330 467 1357 513
rect 1403 467 1440 513
rect 1330 440 1440 467
rect 1380 380 1440 440
rect 1550 380 1610 570
rect 1720 800 1780 1110
rect 1890 930 1950 1110
rect 1890 903 2010 930
rect 1890 857 1937 903
rect 1983 857 2010 903
rect 1890 830 2010 857
rect 1720 773 1840 800
rect 1720 727 1767 773
rect 1813 727 1840 773
rect 1720 700 1840 727
rect 1720 380 1780 700
rect 1890 380 1950 830
rect 2060 540 2120 1110
rect 2230 670 2290 1110
rect 2550 670 2610 1110
rect 2170 643 2290 670
rect 2170 597 2197 643
rect 2243 597 2290 643
rect 2170 570 2290 597
rect 2490 643 2610 670
rect 2490 597 2517 643
rect 2563 597 2610 643
rect 2490 570 2610 597
rect 2010 513 2120 540
rect 2010 467 2037 513
rect 2083 467 2120 513
rect 2010 440 2120 467
rect 2060 380 2120 440
rect 2230 380 2290 570
rect 2550 380 2610 570
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
rect 870 160 930 210
rect 1040 160 1100 210
rect 1210 160 1270 210
rect 1380 160 1440 210
rect 1550 160 1610 210
rect 1720 160 1780 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2550 160 2610 210
<< polycontact >>
rect 327 857 373 903
rect 147 727 193 773
rect 497 597 543 643
rect 747 857 793 903
rect 1177 857 1223 903
rect 947 727 993 773
rect 1517 597 1563 643
rect 1357 467 1403 513
rect 1937 857 1983 903
rect 1767 727 1813 773
rect 2197 597 2243 643
rect 2517 597 2563 643
rect 2037 467 2083 513
<< metal1 >>
rect 0 1588 2800 1670
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1072 1588
rect 1118 1542 1312 1588
rect 1358 1542 1552 1588
rect 1598 1542 1792 1588
rect 1838 1542 2032 1588
rect 2078 1542 2272 1588
rect 2318 1542 2512 1588
rect 2558 1542 2800 1588
rect 0 1520 2800 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1060 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 450 1397 500 1450
rect 450 1163 452 1397
rect 498 1163 500 1397
rect 450 1060 500 1163
rect 110 1010 500 1060
rect 620 1397 670 1450
rect 620 1163 622 1397
rect 668 1163 670 1397
rect 300 906 400 910
rect 300 854 324 906
rect 376 854 400 906
rect 300 850 400 854
rect 120 776 220 780
rect 120 724 144 776
rect 196 724 220 776
rect 120 720 220 724
rect 620 650 670 1163
rect 960 1397 1010 1520
rect 960 1163 962 1397
rect 1008 1163 1010 1397
rect 960 1110 1010 1163
rect 1130 1397 1180 1450
rect 1130 1163 1132 1397
rect 1178 1163 1180 1397
rect 1130 1060 1180 1163
rect 1300 1397 1350 1520
rect 1300 1163 1302 1397
rect 1348 1163 1350 1397
rect 1300 1110 1350 1163
rect 1470 1397 1520 1450
rect 1470 1163 1472 1397
rect 1518 1163 1520 1397
rect 1470 1060 1520 1163
rect 1130 1010 1520 1060
rect 1640 1397 1690 1450
rect 1640 1163 1642 1397
rect 1688 1163 1690 1397
rect 720 906 1250 910
rect 720 854 744 906
rect 796 854 1174 906
rect 1226 854 1250 906
rect 720 850 1250 854
rect 920 776 1020 780
rect 920 724 944 776
rect 996 724 1020 776
rect 920 720 1020 724
rect 1640 650 1690 1163
rect 2150 1397 2200 1520
rect 2150 1163 2152 1397
rect 2198 1163 2200 1397
rect 2150 1110 2200 1163
rect 2320 1397 2370 1450
rect 2320 1163 2322 1397
rect 2368 1163 2370 1397
rect 2320 910 2370 1163
rect 2470 1397 2520 1520
rect 2470 1163 2472 1397
rect 2518 1163 2520 1397
rect 2470 1110 2520 1163
rect 2640 1397 2690 1450
rect 2640 1163 2642 1397
rect 2688 1163 2690 1397
rect 1910 906 2010 910
rect 1910 854 1934 906
rect 1986 854 2010 906
rect 1910 850 2010 854
rect 2320 906 2400 910
rect 2320 854 2324 906
rect 2376 854 2400 906
rect 2320 850 2400 854
rect 1740 776 1840 780
rect 1740 724 1764 776
rect 1816 724 1840 776
rect 1740 720 1840 724
rect 470 646 570 650
rect 470 594 494 646
rect 546 594 570 646
rect 470 590 570 594
rect 620 646 1590 650
rect 620 594 1514 646
rect 1566 594 1590 646
rect 620 590 1590 594
rect 1640 643 2270 650
rect 1640 597 2197 643
rect 2243 597 2270 643
rect 1640 590 2270 597
rect 110 430 500 480
rect 110 318 160 430
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 450 318 500 430
rect 450 272 452 318
rect 498 272 500 318
rect 450 210 500 272
rect 620 318 670 590
rect 1330 516 1430 520
rect 1330 464 1354 516
rect 1406 464 1430 516
rect 1330 460 1430 464
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 960 318 1010 380
rect 960 272 962 318
rect 1008 272 1010 318
rect 960 140 1010 272
rect 1130 360 1520 410
rect 1130 313 1180 360
rect 1130 267 1132 313
rect 1178 267 1180 313
rect 1470 313 1520 360
rect 1130 210 1180 267
rect 1300 283 1350 310
rect 1300 237 1302 283
rect 1348 237 1350 283
rect 1300 140 1350 237
rect 1470 267 1472 313
rect 1518 267 1520 313
rect 1470 210 1520 267
rect 1640 318 1690 590
rect 2010 516 2110 520
rect 2010 464 2034 516
rect 2086 464 2110 516
rect 2010 460 2110 464
rect 1640 272 1642 318
rect 1688 272 1690 318
rect 1640 210 1690 272
rect 2150 318 2200 380
rect 2150 272 2152 318
rect 2198 272 2200 318
rect 2150 140 2200 272
rect 2320 318 2370 850
rect 2640 660 2690 1163
rect 2640 650 2720 660
rect 2490 646 2590 650
rect 2490 594 2514 646
rect 2566 594 2590 646
rect 2490 590 2590 594
rect 2640 646 2750 650
rect 2640 594 2674 646
rect 2726 594 2750 646
rect 2640 590 2750 594
rect 2640 580 2720 590
rect 2320 272 2322 318
rect 2368 272 2370 318
rect 2320 210 2370 272
rect 2470 318 2520 380
rect 2470 272 2472 318
rect 2518 272 2520 318
rect 2470 140 2520 272
rect 2640 318 2690 580
rect 2640 272 2642 318
rect 2688 272 2690 318
rect 2640 210 2690 272
rect 0 118 2800 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2800 118
rect 0 0 2800 72
<< via1 >>
rect 324 903 376 906
rect 324 857 327 903
rect 327 857 373 903
rect 373 857 376 903
rect 324 854 376 857
rect 144 773 196 776
rect 144 727 147 773
rect 147 727 193 773
rect 193 727 196 773
rect 144 724 196 727
rect 744 903 796 906
rect 744 857 747 903
rect 747 857 793 903
rect 793 857 796 903
rect 744 854 796 857
rect 1174 903 1226 906
rect 1174 857 1177 903
rect 1177 857 1223 903
rect 1223 857 1226 903
rect 1174 854 1226 857
rect 944 773 996 776
rect 944 727 947 773
rect 947 727 993 773
rect 993 727 996 773
rect 944 724 996 727
rect 1934 903 1986 906
rect 1934 857 1937 903
rect 1937 857 1983 903
rect 1983 857 1986 903
rect 1934 854 1986 857
rect 2324 854 2376 906
rect 1764 773 1816 776
rect 1764 727 1767 773
rect 1767 727 1813 773
rect 1813 727 1816 773
rect 1764 724 1816 727
rect 494 643 546 646
rect 494 597 497 643
rect 497 597 543 643
rect 543 597 546 643
rect 494 594 546 597
rect 1514 643 1566 646
rect 1514 597 1517 643
rect 1517 597 1563 643
rect 1563 597 1566 643
rect 1514 594 1566 597
rect 1354 513 1406 516
rect 1354 467 1357 513
rect 1357 467 1403 513
rect 1403 467 1406 513
rect 1354 464 1406 467
rect 2034 513 2086 516
rect 2034 467 2037 513
rect 2037 467 2083 513
rect 2083 467 2086 513
rect 2034 464 2086 467
rect 2514 643 2566 646
rect 2514 597 2517 643
rect 2517 597 2563 643
rect 2563 597 2566 643
rect 2514 594 2566 597
rect 2674 594 2726 646
<< metal2 >>
rect 310 910 390 920
rect 730 910 810 920
rect 1160 910 1240 920
rect 1920 910 2000 920
rect 2310 910 2390 920
rect 300 906 820 910
rect 300 854 324 906
rect 376 854 744 906
rect 796 854 820 906
rect 300 850 820 854
rect 1150 906 2010 910
rect 1150 854 1174 906
rect 1226 854 1934 906
rect 1986 854 2010 906
rect 1150 850 2010 854
rect 2300 906 2400 910
rect 2300 854 2324 906
rect 2376 854 2400 906
rect 2300 850 2400 854
rect 310 840 390 850
rect 730 840 810 850
rect 1160 840 1240 850
rect 1920 840 2000 850
rect 2310 840 2390 850
rect 130 780 210 790
rect 930 780 1010 790
rect 1750 780 1830 790
rect 120 776 1840 780
rect 120 724 144 776
rect 196 724 944 776
rect 996 724 1764 776
rect 1816 724 1840 776
rect 120 720 1840 724
rect 130 710 210 720
rect 930 710 1010 720
rect 1750 710 1830 720
rect 480 650 560 660
rect 1500 650 1580 660
rect 2500 650 2580 660
rect 2660 650 2740 660
rect 470 646 570 650
rect 470 594 494 646
rect 546 594 570 646
rect 470 590 570 594
rect 1490 646 2590 650
rect 1490 594 1514 646
rect 1566 594 2514 646
rect 2566 594 2590 646
rect 1490 590 2590 594
rect 2650 646 2750 650
rect 2650 594 2674 646
rect 2726 594 2750 646
rect 2650 590 2750 594
rect 480 580 560 590
rect 1500 580 1580 590
rect 2500 580 2580 590
rect 2660 580 2740 590
rect 490 520 550 580
rect 2510 570 2570 580
rect 1340 520 1420 530
rect 2020 520 2100 530
rect 490 516 2110 520
rect 490 464 1354 516
rect 1406 464 2034 516
rect 2086 464 2110 516
rect 490 460 2110 464
rect 1340 450 1420 460
rect 2020 450 2100 460
rect 1350 440 1410 450
rect 2030 440 2090 450
<< labels >>
rlabel via1 s 1764 724 1816 776 4 A
port 1 nsew signal input
rlabel via1 s 1934 854 1986 906 4 B
port 2 nsew signal input
rlabel via1 s 2034 464 2086 516 4 CI
port 3 nsew signal input
rlabel via1 s 2324 854 2376 906 4 S
port 4 nsew signal output
rlabel via1 s 2674 594 2726 646 4 CO
port 5 nsew signal output
rlabel metal1 s 280 0 330 380 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 280 1110 330 1670 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 960 1110 1010 1670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1300 1110 1350 1670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 1110 2200 1670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2470 1110 2520 1670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1520 2800 1670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 960 0 1010 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1300 0 1350 310 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2150 0 2200 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2470 0 2520 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2800 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel via1 s 944 724 996 776 1 A
port 1 nsew signal input
rlabel via1 s 144 724 196 776 1 A
port 1 nsew signal input
rlabel metal2 s 130 710 210 790 1 A
port 1 nsew signal input
rlabel metal2 s 930 710 1010 790 1 A
port 1 nsew signal input
rlabel metal2 s 1750 710 1830 790 1 A
port 1 nsew signal input
rlabel metal2 s 120 720 1840 780 1 A
port 1 nsew signal input
rlabel metal1 s 120 720 220 780 1 A
port 1 nsew signal input
rlabel metal1 s 920 720 1020 780 1 A
port 1 nsew signal input
rlabel metal1 s 1740 720 1840 780 1 A
port 1 nsew signal input
rlabel via1 s 1174 854 1226 906 1 B
port 2 nsew signal input
rlabel via1 s 744 854 796 906 1 B
port 2 nsew signal input
rlabel via1 s 324 854 376 906 1 B
port 2 nsew signal input
rlabel metal2 s 310 840 390 920 1 B
port 2 nsew signal input
rlabel metal2 s 730 840 810 920 1 B
port 2 nsew signal input
rlabel metal2 s 300 850 820 910 1 B
port 2 nsew signal input
rlabel metal2 s 1160 840 1240 920 1 B
port 2 nsew signal input
rlabel metal2 s 1920 840 2000 920 1 B
port 2 nsew signal input
rlabel metal2 s 1150 850 2010 910 1 B
port 2 nsew signal input
rlabel metal1 s 300 850 400 910 1 B
port 2 nsew signal input
rlabel metal1 s 720 850 1250 910 1 B
port 2 nsew signal input
rlabel metal1 s 1910 850 2010 910 1 B
port 2 nsew signal input
rlabel via1 s 1354 464 1406 516 1 CI
port 3 nsew signal input
rlabel via1 s 494 594 546 646 1 CI
port 3 nsew signal input
rlabel metal2 s 490 460 550 660 1 CI
port 3 nsew signal input
rlabel metal2 s 480 580 560 660 1 CI
port 3 nsew signal input
rlabel metal2 s 470 590 570 650 1 CI
port 3 nsew signal input
rlabel metal2 s 1350 440 1410 530 1 CI
port 3 nsew signal input
rlabel metal2 s 1340 450 1420 530 1 CI
port 3 nsew signal input
rlabel metal2 s 2030 440 2090 530 1 CI
port 3 nsew signal input
rlabel metal2 s 2020 450 2100 530 1 CI
port 3 nsew signal input
rlabel metal2 s 490 460 2110 520 1 CI
port 3 nsew signal input
rlabel metal1 s 470 590 570 650 1 CI
port 3 nsew signal input
rlabel metal1 s 1330 460 1430 520 1 CI
port 3 nsew signal input
rlabel metal1 s 2010 460 2110 520 1 CI
port 3 nsew signal input
rlabel metal2 s 2660 580 2740 660 1 CO
port 5 nsew signal output
rlabel metal2 s 2650 590 2750 650 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 210 2690 1450 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 580 2720 660 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 590 2750 650 1 CO
port 5 nsew signal output
rlabel metal2 s 2310 840 2390 920 1 S
port 4 nsew signal output
rlabel metal2 s 2300 850 2400 910 1 S
port 4 nsew signal output
rlabel metal1 s 2320 210 2370 1450 1 S
port 4 nsew signal output
rlabel metal1 s 2320 850 2400 910 1 S
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2800 1670
string GDS_END 19172
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 146
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
