magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 982 1094
<< pwell >>
rect -86 -86 982 453
<< metal1 >>
rect 0 918 896 1098
rect 69 710 115 918
rect 142 443 203 542
rect 360 454 428 542
rect 590 354 642 511
rect 701 296 767 872
rect 273 250 767 296
rect 49 90 95 204
rect 273 136 319 250
rect 497 90 543 204
rect 721 136 767 250
rect 0 -90 896 90
<< labels >>
rlabel metal1 s 590 354 642 511 6 A1
port 1 nsew default input
rlabel metal1 s 360 454 428 542 6 A2
port 2 nsew default input
rlabel metal1 s 142 443 203 542 6 A3
port 3 nsew default input
rlabel metal1 s 721 136 767 250 6 ZN
port 4 nsew default output
rlabel metal1 s 273 136 319 250 6 ZN
port 4 nsew default output
rlabel metal1 s 273 250 767 296 6 ZN
port 4 nsew default output
rlabel metal1 s 701 296 767 872 6 ZN
port 4 nsew default output
rlabel metal1 s 69 710 115 918 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 918 896 1098 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 453 982 1094 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 982 453 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -90 896 90 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 204 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 204 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 88632
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 85734
<< end >>
