VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__dvss
  CLASS PAD POWER ;
  FOREIGN gf180mcu_fd_io__dvss ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 62.490 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.490 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 12.510 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 12.510 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 12.510 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 12.510 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 12.510 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 12.510 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 12.510 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 12.510 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 12.510 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 12.510 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 12.510 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 12.510 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 1.360 349.000 10.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 13.760 349.000 24.010 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 25.610 349.000 35.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 39.140 349.000 49.390 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 50.990 349.000 61.240 350.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 64.140 349.000 73.640 350.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 11.845 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.845 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 11.565 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 11.565 261.000 ;
    END
  END VDD
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 348.700 1.060 349.000 ;
        RECT 11.160 348.700 13.460 349.000 ;
        RECT 24.310 348.700 25.310 349.000 ;
        RECT 36.160 348.700 38.840 349.000 ;
        RECT 49.690 348.700 50.690 349.000 ;
        RECT 61.540 348.700 63.840 349.000 ;
        RECT 73.940 348.700 75.000 349.000 ;
        RECT 0.000 0.000 75.000 348.700 ;
      LAYER Metal3 ;
        RECT 2.800 342.800 72.200 348.390 ;
        RECT 14.310 332.200 60.690 342.800 ;
        RECT 2.800 318.800 72.200 332.200 ;
        RECT 2.800 302.800 72.200 308.200 ;
        RECT 14.310 292.200 60.690 302.800 ;
        RECT 2.800 286.800 72.200 292.200 ;
        RECT 14.310 262.800 60.690 286.800 ;
        RECT 2.800 230.800 72.200 252.200 ;
        RECT 14.310 204.200 60.690 230.800 ;
        RECT 2.800 198.800 72.200 204.200 ;
        RECT 14.310 132.200 60.690 198.800 ;
        RECT 2.800 126.800 72.200 132.200 ;
        RECT 14.310 116.200 60.690 126.800 ;
        RECT 2.800 68.200 72.200 116.200 ;
        RECT 1.000 0.000 74.000 68.200 ;
  END
END gf180mcu_fd_io__dvss
END LIBRARY

