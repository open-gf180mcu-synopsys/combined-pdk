magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1070 1270
<< nmos >>
rect 190 210 250 380
rect 380 210 440 380
rect 490 210 550 380
rect 810 210 870 380
<< pmos >>
rect 190 720 250 1060
rect 380 720 440 1060
rect 490 720 550 1060
rect 810 720 870 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 380 380
rect 250 272 292 318
rect 338 272 380 318
rect 250 210 380 272
rect 440 210 490 380
rect 550 318 650 380
rect 550 272 582 318
rect 628 272 650 318
rect 550 210 650 272
rect 710 318 810 380
rect 710 272 732 318
rect 778 272 810 318
rect 710 210 810 272
rect 870 318 970 380
rect 870 272 902 318
rect 948 272 970 318
rect 870 210 970 272
<< pdiff >>
rect 90 1000 190 1060
rect 90 860 112 1000
rect 158 860 190 1000
rect 90 720 190 860
rect 250 1000 380 1060
rect 250 860 292 1000
rect 338 860 380 1000
rect 250 720 380 860
rect 440 720 490 1060
rect 550 1007 650 1060
rect 550 773 582 1007
rect 628 773 650 1007
rect 550 720 650 773
rect 710 1007 810 1060
rect 710 773 732 1007
rect 778 773 810 1007
rect 710 720 810 773
rect 870 1005 970 1060
rect 870 865 902 1005
rect 948 865 970 1005
rect 870 720 970 865
<< ndiffc >>
rect 112 272 158 318
rect 292 272 338 318
rect 582 272 628 318
rect 732 272 778 318
rect 902 272 948 318
<< pdiffc >>
rect 112 860 158 1000
rect 292 860 338 1000
rect 582 773 628 1007
rect 732 773 778 1007
rect 902 865 948 1005
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 290 1198 440 1220
rect 290 1152 342 1198
rect 388 1152 440 1198
rect 290 1130 440 1152
rect 520 1198 670 1220
rect 520 1152 572 1198
rect 618 1152 670 1198
rect 520 1130 670 1152
rect 750 1198 900 1220
rect 750 1152 802 1198
rect 848 1152 900 1198
rect 750 1130 900 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 342 1152 388 1198
rect 572 1152 618 1198
rect 802 1152 848 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 380 1060 440 1110
rect 490 1060 550 1110
rect 810 1060 870 1110
rect 190 670 250 720
rect 190 643 290 670
rect 190 597 217 643
rect 263 597 290 643
rect 190 570 290 597
rect 190 380 250 570
rect 380 520 440 720
rect 490 640 550 720
rect 610 640 710 660
rect 490 638 710 640
rect 490 592 642 638
rect 688 592 710 638
rect 490 580 710 592
rect 610 570 710 580
rect 810 530 870 720
rect 750 520 870 530
rect 330 493 440 520
rect 330 447 357 493
rect 403 447 440 493
rect 330 420 440 447
rect 380 380 440 420
rect 490 508 870 520
rect 490 462 782 508
rect 828 462 870 508
rect 490 460 870 462
rect 490 380 550 460
rect 750 440 870 460
rect 810 380 870 440
rect 190 160 250 210
rect 380 160 440 210
rect 490 160 550 210
rect 810 160 870 210
<< polycontact >>
rect 217 597 263 643
rect 642 592 688 638
rect 357 447 403 493
rect 782 462 828 508
<< metal1 >>
rect 0 1198 1070 1270
rect 0 1152 112 1198
rect 158 1152 342 1198
rect 388 1152 572 1198
rect 618 1152 802 1198
rect 848 1152 1070 1198
rect 0 1130 1070 1152
rect 110 1000 160 1060
rect 110 860 112 1000
rect 158 860 160 1000
rect 110 780 160 860
rect 280 1000 350 1130
rect 280 860 292 1000
rect 338 860 350 1000
rect 280 800 350 860
rect 580 1007 630 1060
rect 90 700 160 780
rect 580 773 582 1007
rect 628 930 630 1007
rect 730 1007 780 1130
rect 628 906 640 930
rect 636 854 640 906
rect 628 830 640 854
rect 628 773 630 830
rect 580 750 630 773
rect 490 700 630 750
rect 730 773 732 1007
rect 778 773 780 1007
rect 730 720 780 773
rect 900 1005 950 1060
rect 900 865 902 1005
rect 948 865 950 1005
rect 90 500 140 700
rect 190 646 290 650
rect 190 594 214 646
rect 266 594 290 646
rect 190 590 290 594
rect 90 493 430 500
rect 90 447 357 493
rect 403 447 430 493
rect 90 440 430 447
rect 90 380 140 440
rect 490 380 540 700
rect 900 650 950 865
rect 610 646 950 650
rect 610 594 634 646
rect 686 638 950 646
rect 610 592 642 594
rect 688 592 950 638
rect 610 590 950 592
rect 750 516 850 520
rect 750 464 774 516
rect 826 508 850 516
rect 750 462 782 464
rect 828 462 850 508
rect 750 460 850 462
rect 90 320 160 380
rect 110 318 160 320
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 350 380
rect 490 330 630 380
rect 280 272 292 318
rect 338 272 350 318
rect 280 140 350 272
rect 580 318 630 330
rect 580 272 582 318
rect 628 272 630 318
rect 580 210 630 272
rect 730 318 780 380
rect 730 272 732 318
rect 778 272 780 318
rect 730 140 780 272
rect 900 318 950 590
rect 900 272 902 318
rect 948 272 950 318
rect 900 210 950 272
rect 0 118 1070 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1070 118
rect 0 0 1070 72
<< via1 >>
rect 584 854 628 906
rect 628 854 636 906
rect 214 643 266 646
rect 214 597 217 643
rect 217 597 263 643
rect 263 597 266 643
rect 214 594 266 597
rect 634 638 686 646
rect 634 594 642 638
rect 642 594 686 638
rect 774 508 826 516
rect 774 464 782 508
rect 782 464 826 508
<< metal2 >>
rect 560 906 660 920
rect 560 854 584 906
rect 636 854 660 906
rect 560 840 660 854
rect 200 650 280 660
rect 190 646 290 650
rect 190 594 214 646
rect 266 594 290 646
rect 190 590 290 594
rect 610 646 710 660
rect 610 594 634 646
rect 686 594 710 646
rect 200 580 280 590
rect 610 580 710 594
rect 750 516 850 530
rect 750 464 774 516
rect 826 464 850 516
rect 750 450 850 464
<< labels >>
rlabel via1 s 214 594 266 646 4 A
port 1 nsew signal input
rlabel via1 s 584 854 636 906 4 Y
port 2 nsew signal output
rlabel via1 s 774 464 826 516 4 EN
port 3 nsew signal input
rlabel metal1 s 280 800 350 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 350 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 730 720 780 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1070 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 730 0 780 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1070 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 200 580 280 660 1 A
port 1 nsew signal input
rlabel metal2 s 190 590 290 650 1 A
port 1 nsew signal input
rlabel metal1 s 190 590 290 650 1 A
port 1 nsew signal input
rlabel metal2 s 750 450 850 530 1 EN
port 3 nsew signal input
rlabel metal1 s 750 460 850 520 1 EN
port 3 nsew signal input
rlabel metal2 s 560 840 660 920 1 Y
port 2 nsew signal output
rlabel metal1 s 490 330 540 750 1 Y
port 2 nsew signal output
rlabel metal1 s 490 700 630 750 1 Y
port 2 nsew signal output
rlabel metal1 s 580 210 630 380 1 Y
port 2 nsew signal output
rlabel metal1 s 490 330 630 380 1 Y
port 2 nsew signal output
rlabel metal1 s 580 700 630 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 580 830 640 930 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1070 1270
string GDS_END 367416
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 360498
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
