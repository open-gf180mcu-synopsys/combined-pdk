magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 3110 1094
<< pwell >>
rect -86 -86 3110 453
<< mvnmos >>
rect 168 156 288 296
rect 392 156 512 296
rect 616 156 736 296
rect 840 156 960 296
rect 1008 156 1128 296
rect 1232 156 1352 296
rect 1703 137 1823 277
rect 1927 137 2047 277
rect 2295 137 2415 277
rect 2463 137 2583 277
rect 2727 133 2847 333
<< mvpmos >>
rect 244 576 344 852
rect 392 576 492 852
rect 544 576 644 852
rect 928 576 1028 852
rect 1076 576 1176 852
rect 1280 576 1380 852
rect 1713 577 1813 853
rect 1917 577 2017 853
rect 2269 573 2369 849
rect 2473 573 2573 849
rect 2713 573 2813 939
<< mvndiff >>
rect 36 196 168 296
rect 36 150 49 196
rect 95 156 168 196
rect 288 215 392 296
rect 288 169 317 215
rect 363 169 392 215
rect 288 156 392 169
rect 512 215 616 296
rect 512 169 541 215
rect 587 169 616 215
rect 512 156 616 169
rect 736 215 840 296
rect 736 169 765 215
rect 811 169 840 215
rect 736 156 840 169
rect 960 156 1008 296
rect 1128 215 1232 296
rect 1128 169 1157 215
rect 1203 169 1232 215
rect 1128 156 1232 169
rect 1352 215 1440 296
rect 1352 169 1381 215
rect 1427 169 1440 215
rect 1352 156 1440 169
rect 95 150 108 156
rect 36 137 108 150
rect 2647 277 2727 333
rect 1615 196 1703 277
rect 1615 150 1628 196
rect 1674 150 1703 196
rect 1615 137 1703 150
rect 1823 196 1927 277
rect 1823 150 1852 196
rect 1898 150 1927 196
rect 1823 137 1927 150
rect 2047 196 2135 277
rect 2047 150 2076 196
rect 2122 150 2135 196
rect 2047 137 2135 150
rect 2207 196 2295 277
rect 2207 150 2220 196
rect 2266 150 2295 196
rect 2207 137 2295 150
rect 2415 137 2463 277
rect 2583 192 2727 277
rect 2583 146 2652 192
rect 2698 146 2727 192
rect 2583 137 2727 146
rect 2643 133 2727 137
rect 2847 290 2935 333
rect 2847 150 2876 290
rect 2922 150 2935 290
rect 2847 133 2935 150
<< mvpdiff >>
rect 156 838 244 852
rect 156 698 169 838
rect 215 698 244 838
rect 156 576 244 698
rect 344 576 392 852
rect 492 576 544 852
rect 644 838 928 852
rect 644 698 673 838
rect 719 698 928 838
rect 644 576 928 698
rect 1028 576 1076 852
rect 1176 839 1280 852
rect 1176 793 1205 839
rect 1251 793 1280 839
rect 1176 576 1280 793
rect 1380 838 1468 852
rect 1380 698 1409 838
rect 1455 698 1468 838
rect 1380 576 1468 698
rect 1625 636 1713 853
rect 1625 590 1638 636
rect 1684 590 1713 636
rect 1625 577 1713 590
rect 1813 836 1917 853
rect 1813 790 1842 836
rect 1888 790 1917 836
rect 1813 577 1917 790
rect 2017 636 2105 853
rect 2633 849 2713 939
rect 2017 590 2046 636
rect 2092 590 2105 636
rect 2017 577 2105 590
rect 2181 836 2269 849
rect 2181 790 2194 836
rect 2240 790 2269 836
rect 2181 573 2269 790
rect 2369 726 2473 849
rect 2369 586 2398 726
rect 2444 586 2473 726
rect 2369 573 2473 586
rect 2573 836 2713 849
rect 2573 696 2602 836
rect 2648 696 2713 836
rect 2573 573 2713 696
rect 2813 726 2901 939
rect 2813 586 2842 726
rect 2888 586 2901 726
rect 2813 573 2901 586
<< mvndiffc >>
rect 49 150 95 196
rect 317 169 363 215
rect 541 169 587 215
rect 765 169 811 215
rect 1157 169 1203 215
rect 1381 169 1427 215
rect 1628 150 1674 196
rect 1852 150 1898 196
rect 2076 150 2122 196
rect 2220 150 2266 196
rect 2652 146 2698 192
rect 2876 150 2922 290
<< mvpdiffc >>
rect 169 698 215 838
rect 673 698 719 838
rect 1205 793 1251 839
rect 1409 698 1455 838
rect 1638 590 1684 636
rect 1842 790 1888 836
rect 2046 590 2092 636
rect 2194 790 2240 836
rect 2398 586 2444 726
rect 2602 696 2648 836
rect 2842 586 2888 726
<< polysilicon >>
rect 928 944 1813 984
rect 244 852 344 896
rect 392 852 492 896
rect 544 852 644 896
rect 928 852 1028 944
rect 1076 852 1176 896
rect 1280 852 1380 896
rect 1713 853 1813 944
rect 2713 939 2813 983
rect 1917 853 2017 897
rect 2269 849 2369 893
rect 2473 849 2573 893
rect 244 532 344 576
rect 244 513 288 532
rect 168 500 288 513
rect 168 454 181 500
rect 227 454 288 500
rect 168 296 288 454
rect 392 500 492 576
rect 392 454 405 500
rect 451 454 492 500
rect 544 516 644 576
rect 928 543 1028 576
rect 544 476 880 516
rect 928 497 941 543
rect 987 497 1028 543
rect 928 484 1028 497
rect 1076 513 1176 576
rect 1280 532 1380 576
rect 1076 500 1195 513
rect 392 340 492 454
rect 616 415 792 428
rect 616 369 733 415
rect 779 369 792 415
rect 616 356 792 369
rect 392 296 512 340
rect 616 296 736 356
rect 840 340 880 476
rect 1076 454 1136 500
rect 1182 454 1195 500
rect 1076 441 1195 454
rect 1280 500 1352 532
rect 1280 454 1293 500
rect 1339 454 1352 500
rect 1076 340 1128 441
rect 1280 340 1352 454
rect 840 296 960 340
rect 1008 296 1128 340
rect 1232 296 1352 340
rect 1511 521 1583 534
rect 1511 475 1524 521
rect 1570 475 1583 521
rect 1511 462 1583 475
rect 1713 500 1813 577
rect 168 112 288 156
rect 392 112 512 156
rect 616 112 736 156
rect 840 64 960 156
rect 1008 112 1128 156
rect 1232 112 1352 156
rect 1511 64 1551 462
rect 1713 454 1754 500
rect 1800 454 1813 500
rect 1713 321 1813 454
rect 1917 513 2017 577
rect 2269 513 2369 573
rect 2473 513 2573 573
rect 1917 500 2369 513
rect 1917 454 2046 500
rect 2092 454 2369 500
rect 1917 441 2369 454
rect 2441 500 2573 513
rect 2441 454 2454 500
rect 2500 454 2573 500
rect 2441 441 2573 454
rect 2713 500 2813 573
rect 2713 454 2726 500
rect 2772 454 2813 500
rect 2713 441 2813 454
rect 1917 359 2047 441
rect 1703 277 1823 321
rect 1927 277 2047 359
rect 2295 321 2369 441
rect 2463 321 2573 441
rect 2727 377 2813 441
rect 2727 333 2847 377
rect 2295 277 2415 321
rect 2463 277 2583 321
rect 1703 93 1823 137
rect 1927 93 2047 137
rect 2295 93 2415 137
rect 2463 93 2583 137
rect 2727 89 2847 133
rect 840 24 1551 64
<< polycontact >>
rect 181 454 227 500
rect 405 454 451 500
rect 941 497 987 543
rect 733 369 779 415
rect 1136 454 1182 500
rect 1293 454 1339 500
rect 1524 475 1570 521
rect 1754 454 1800 500
rect 2046 454 2092 500
rect 2454 454 2500 500
rect 2726 454 2772 500
<< metal1 >>
rect 0 918 3024 1098
rect 169 838 215 918
rect 169 687 215 698
rect 641 838 719 849
rect 641 698 673 838
rect 1205 839 1251 918
rect 1205 782 1251 793
rect 1409 838 1455 849
rect 641 635 719 698
rect 1136 698 1409 728
rect 1796 847 1842 918
rect 1796 836 2648 847
rect 1796 790 1842 836
rect 1888 790 2194 836
rect 2240 801 2602 836
rect 1796 779 2240 790
rect 1455 698 2195 728
rect 1136 682 2195 698
rect 641 589 1090 635
rect 366 500 451 542
rect 30 454 181 500
rect 227 454 238 500
rect 366 454 405 500
rect 30 242 82 454
rect 366 354 451 454
rect 128 261 587 307
rect 128 196 174 261
rect 541 215 587 261
rect 38 150 49 196
rect 95 150 174 196
rect 306 169 317 215
rect 363 169 374 215
rect 306 90 374 169
rect 641 215 687 589
rect 733 497 941 543
rect 987 497 998 543
rect 733 415 779 497
rect 733 358 779 369
rect 1044 397 1090 589
rect 1136 500 1182 682
rect 1136 443 1182 454
rect 1228 454 1293 500
rect 1339 454 1350 500
rect 1228 397 1274 454
rect 1044 351 1274 397
rect 1396 226 1442 682
rect 1627 590 1638 636
rect 1684 590 1695 636
rect 1627 521 1695 590
rect 1513 475 1524 521
rect 1570 475 1695 521
rect 1954 590 2046 636
rect 2092 590 2103 636
rect 1954 500 2000 590
rect 1157 215 1203 226
rect 641 169 765 215
rect 811 169 822 215
rect 541 158 587 169
rect 1157 90 1203 169
rect 1381 215 1442 226
rect 1427 169 1442 215
rect 1381 158 1442 169
rect 1628 196 1695 475
rect 1743 454 1754 500
rect 1800 454 2000 500
rect 1674 150 1695 196
rect 1628 139 1695 150
rect 1852 196 1898 207
rect 1954 196 2000 454
rect 2046 500 2098 542
rect 2092 454 2098 500
rect 2149 500 2195 682
rect 2398 726 2444 737
rect 2602 685 2648 696
rect 2830 726 2922 737
rect 2444 586 2603 621
rect 2398 575 2603 586
rect 2557 500 2603 575
rect 2830 586 2842 726
rect 2888 586 2922 726
rect 2149 454 2454 500
rect 2500 454 2511 500
rect 2557 454 2726 500
rect 2772 454 2783 500
rect 2046 354 2098 454
rect 2557 207 2603 454
rect 2220 196 2603 207
rect 2830 290 2922 586
rect 1954 150 2076 196
rect 2122 150 2133 196
rect 2266 150 2603 196
rect 1852 90 1898 150
rect 2220 139 2603 150
rect 2652 192 2698 203
rect 2652 90 2698 146
rect 2830 150 2876 290
rect 2830 139 2922 150
rect 0 -90 3024 90
<< labels >>
flabel metal1 s 2046 354 2098 542 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 366 354 451 542 0 FreeSans 200 0 0 0 E
port 2 nsew default input
flabel metal1 s 2830 139 2922 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 30 454 238 500 0 FreeSans 200 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 918 3024 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1157 215 1203 226 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 30 242 82 454 1 TE
port 3 nsew default input
rlabel metal1 s 1796 847 1842 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1205 847 1251 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 169 847 215 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1796 801 2648 847 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1205 801 1251 847 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 169 801 215 847 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2602 782 2648 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1796 782 2240 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1205 782 1251 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 169 782 215 801 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2602 779 2648 782 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1796 779 2240 782 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 169 779 215 782 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2602 687 2648 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 169 687 215 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2602 685 2648 687 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1157 207 1203 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 306 207 374 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1852 203 1898 207 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1157 203 1203 207 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 306 203 374 207 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2652 90 2698 203 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1852 90 1898 203 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1157 90 1203 203 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 306 90 374 203 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3024 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3024 1008
string GDS_END 852380
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 845304
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
