magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use M1_NWELL$$47634476_64x8m81  M1_NWELL$$47634476_64x8m81_0
timestamp 1750858719
transform 1 0 9487 0 1 16304
box 0 0 1 1
use M1_NWELL$$47635500_64x8m81  M1_NWELL$$47635500_64x8m81_0
timestamp 1750858719
transform 1 0 10211 0 1 442
box 0 0 1 1
use M1_POLY24310589983234_64x8m81  M1_POLY24310589983234_64x8m81_0
timestamp 1750858719
transform 1 0 6424 0 1 179
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1750858719
transform 1 0 7216 0 1 849
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1750858719
transform 0 -1 8151 1 0 865
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_1
timestamp 1750858719
transform 1 0 7471 0 1 1141
box 0 0 1 1
use M1_PSUB$$47114284_64x8m81  M1_PSUB$$47114284_64x8m81_0
timestamp 1750858719
transform 1 0 10240 0 1 1283
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1750858719
transform -1 0 7466 0 1 1231
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1750858719
transform -1 0 5683 0 1 732
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_2
timestamp 1750858719
transform -1 0 6303 0 1 1181
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_3
timestamp 1750858719
transform -1 0 6939 0 1 483
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_4
timestamp 1750858719
transform -1 0 5912 0 1 465
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_0
timestamp 1750858719
transform -1 0 5202 0 1 3546
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_1
timestamp 1750858719
transform -1 0 4688 0 1 4151
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_2
timestamp 1750858719
transform -1 0 1820 0 1 3949
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_3
timestamp 1750858719
transform -1 0 3511 0 1 3747
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_4
timestamp 1750858719
transform -1 0 2998 0 1 4353
box 0 0 1 1
use M2_M1$$47630380_64x8m81  M2_M1$$47630380_64x8m81_0
timestamp 1750858719
transform -1 0 10023 0 1 478
box 0 0 1 1
use M2_M1$$47631404_64x8m81  M2_M1$$47631404_64x8m81_0
timestamp 1750858719
transform -1 0 10157 0 1 1313
box 0 0 1 1
use M2_M14310589983217_64x8m81  M2_M14310589983217_64x8m81_0
timestamp 1750858719
transform 1 0 7211 0 1 865
box 0 0 1 1
use M2_M14310589983217_64x8m81  M2_M14310589983217_64x8m81_1
timestamp 1750858719
transform 1 0 8182 0 1 865
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_0
timestamp 1750858719
transform -1 0 6303 0 1 1181
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_1
timestamp 1750858719
transform -1 0 6939 0 1 483
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_2
timestamp 1750858719
transform -1 0 5912 0 1 465
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_3
timestamp 1750858719
transform 1 0 2712 0 1 10925
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_4
timestamp 1750858719
transform 1 0 472 0 1 11455
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_5
timestamp 1750858719
transform 1 0 11208 0 1 11471
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_6
timestamp 1750858719
transform 1 0 12792 0 1 10975
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_7
timestamp 1750858719
transform 1 0 13912 0 1 10766
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_8
timestamp 1750858719
transform 1 0 15032 0 1 10557
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_9
timestamp 1750858719
transform 1 0 16152 0 1 10349
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_10
timestamp 1750858719
transform 1 0 17272 0 1 10140
box 0 0 1 1
use M3_M2$$43368492_R90_64x8m81  M3_M2$$43368492_R90_64x8m81_0
timestamp 1750858719
transform 0 -1 10657 1 0 11262
box 0 0 1 1
use M3_M2$$43368492_R270_64x8m81  M3_M2$$43368492_R270_64x8m81_0
timestamp 1750858719
transform 0 1 11777 -1 0 11061
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_0
timestamp 1750858719
transform 1 0 8841 0 1 10637
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_1
timestamp 1750858719
transform 1 0 6999 0 1 10220
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_2
timestamp 1750858719
transform 1 0 6362 0 1 10011
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_3
timestamp 1750858719
transform 1 0 8417 0 1 10011
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_4
timestamp 1750858719
transform 1 0 7890 0 1 10428
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_5
timestamp 1750858719
transform 1 0 6072 0 1 10428
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_6
timestamp 1750858719
transform 1 0 4952 0 1 10637
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_7
timestamp 1750858719
transform 1 0 3937 0 1 10845
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_8
timestamp 1750858719
transform 1 0 1698 0 1 11262
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_9
timestamp 1750858719
transform 1 0 9524 0 1 10845
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_10
timestamp 1750858719
transform 1 0 9537 0 1 11471
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_0
timestamp 1750858719
transform 1 0 6953 0 1 13665
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_1
timestamp 1750858719
transform 1 0 6505 0 1 13665
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_2
timestamp 1750858719
transform 1 0 8072 0 1 14006
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_3
timestamp 1750858719
transform 1 0 7625 0 1 14006
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_4
timestamp 1750858719
transform 1 0 9192 0 1 14346
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_5
timestamp 1750858719
transform 1 0 8744 0 1 14346
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_6
timestamp 1750858719
transform 1 0 905 0 1 11965
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_7
timestamp 1750858719
transform 1 0 1353 0 1 11965
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_8
timestamp 1750858719
transform 1 0 2473 0 1 12305
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_9
timestamp 1750858719
transform 1 0 2025 0 1 12305
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_10
timestamp 1750858719
transform 1 0 3593 0 1 12645
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_11
timestamp 1750858719
transform 1 0 3145 0 1 12645
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_12
timestamp 1750858719
transform 1 0 4713 0 1 12985
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_13
timestamp 1750858719
transform 1 0 4265 0 1 12985
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_14
timestamp 1750858719
transform 1 0 5833 0 1 13325
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_15
timestamp 1750858719
transform 1 0 5385 0 1 13325
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_16
timestamp 1750858719
transform -1 0 11432 0 -1 12305
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_17
timestamp 1750858719
transform -1 0 10984 0 -1 12305
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_18
timestamp 1750858719
transform -1 0 12552 0 -1 12645
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_19
timestamp 1750858719
transform -1 0 12104 0 -1 12645
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_20
timestamp 1750858719
transform -1 0 13672 0 -1 12985
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_21
timestamp 1750858719
transform -1 0 13224 0 -1 12985
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_22
timestamp 1750858719
transform -1 0 14792 0 -1 13325
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_23
timestamp 1750858719
transform -1 0 14344 0 -1 13325
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_24
timestamp 1750858719
transform -1 0 15912 0 -1 13665
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_25
timestamp 1750858719
transform -1 0 15464 0 -1 13665
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_26
timestamp 1750858719
transform -1 0 17032 0 -1 14006
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_27
timestamp 1750858719
transform -1 0 16584 0 -1 14006
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_28
timestamp 1750858719
transform -1 0 17704 0 -1 14346
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_29
timestamp 1750858719
transform -1 0 18152 0 -1 14346
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_30
timestamp 1750858719
transform 1 0 10086 0 1 11054
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_31
timestamp 1750858719
transform -1 0 10312 0 -1 11965
box 0 0 1 1
use M3_M2$$46895148_64x8m81  M3_M2$$46895148_64x8m81_32
timestamp 1750858719
transform -1 0 9864 0 -1 11965
box 0 0 1 1
use M3_M2$$47632428_64x8m81  M3_M2$$47632428_64x8m81_0
timestamp 1750858719
transform -1 0 10023 0 1 478
box 0 0 1 1
use M3_M2$$47633452_64x8m81  M3_M2$$47633452_64x8m81_0
timestamp 1750858719
transform -1 0 10157 0 1 1313
box 0 0 1 1
use nmos_1p2$$47342636_64x8m81  nmos_1p2$$47342636_64x8m81_0
timestamp 1750858719
transform -1 0 6441 0 1 997
box -31 0 -30 1
use nmos_5p04310589983260_64x8m81  nmos_5p04310589983260_64x8m81_0
timestamp 1750858719
transform -1 0 7842 0 1 1002
box 0 0 1 1
use nmos_5p04310589983260_64x8m81  nmos_5p04310589983260_64x8m81_1
timestamp 1750858719
transform -1 0 8066 0 1 1002
box 0 0 1 1
use pmos_1p2$$47109164_64x8m81  pmos_1p2$$47109164_64x8m81_0
timestamp 1750858719
transform -1 0 6559 0 1 281
box -31 0 -30 1
use ypredec1_bot_64x8m81  ypredec1_bot_64x8m81_0
timestamp 1750858719
transform 1 0 3766 0 1 1027
box -20 -633 1762 7425
use ypredec1_bot_64x8m81  ypredec1_bot_64x8m81_1
timestamp 1750858719
transform 1 0 384 0 1 1027
box -20 -633 1762 7425
use ypredec1_bot_64x8m81  ypredec1_bot_64x8m81_2
timestamp 1750858719
transform 1 0 2075 0 1 1027
box -20 -633 1762 7425
use ypredec1_xax8_64x8m81  ypredec1_xax8_64x8m81_0
timestamp 1750858719
transform 1 0 5624 0 1 1528
box 287 1002 6534 6933
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_0
timestamp 1750858719
transform 1 0 255 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_1
timestamp 1750858719
transform 1 0 1375 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_2
timestamp 1750858719
transform 1 0 2495 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_3
timestamp 1750858719
transform 1 0 3615 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_4
timestamp 1750858719
transform 1 0 4735 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_5
timestamp 1750858719
transform 1 0 5855 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_6
timestamp 1750858719
transform 1 0 6975 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_7
timestamp 1750858719
transform 1 0 10335 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_8
timestamp 1750858719
transform 1 0 11455 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_9
timestamp 1750858719
transform 1 0 12575 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_10
timestamp 1750858719
transform 1 0 13695 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_11
timestamp 1750858719
transform 1 0 14815 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_12
timestamp 1750858719
transform 1 0 15935 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_13
timestamp 1750858719
transform 1 0 17055 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_14
timestamp 1750858719
transform 1 0 9215 0 1 9054
box 202 340 1323 6581
use ypredec1_ys_64x8m81  ypredec1_ys_64x8m81_15
timestamp 1750858719
transform 1 0 8095 0 1 9054
box 202 340 1323 6581
<< properties >>
string GDS_END 1436748
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1415262
<< end >>
