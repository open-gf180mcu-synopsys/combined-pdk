magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< psubdiff >>
rect 0 69946 400 69968
rect 0 69897 127 69946
rect 273 69897 400 69946
rect 0 13151 25 69897
rect 71 69778 329 69800
rect 71 13287 93 69778
rect 307 13287 329 69778
rect 71 13265 329 13287
rect 375 13151 400 69897
rect 0 13119 127 13151
rect 273 13119 400 13151
rect 0 13097 400 13119
<< psubdiffcont >>
rect 127 69897 273 69946
rect 25 69800 375 69897
rect 25 13265 71 69800
rect 329 13265 375 69800
rect 25 13151 375 13265
rect 127 13119 273 13151
<< metal1 >>
rect -32 69946 432 69957
rect -32 69897 127 69946
rect 273 69897 432 69946
rect -32 13151 25 69897
rect 71 69789 329 69800
rect 71 64990 82 69789
rect 318 64990 329 69789
rect 71 64942 329 64990
rect 71 64890 130 64942
rect 286 64890 329 64942
rect 71 64830 329 64890
rect 71 64778 130 64830
rect 286 64778 329 64830
rect 71 64718 329 64778
rect 71 64666 130 64718
rect 286 64666 329 64718
rect 71 64606 329 64666
rect 71 64554 130 64606
rect 286 64554 329 64606
rect 71 64494 329 64554
rect 71 64442 130 64494
rect 286 64442 329 64494
rect 71 64382 329 64442
rect 71 64330 130 64382
rect 286 64330 329 64382
rect 71 64270 329 64330
rect 71 64218 130 64270
rect 286 64218 329 64270
rect 71 64158 329 64218
rect 71 64106 130 64158
rect 286 64106 329 64158
rect 71 64046 329 64106
rect 71 63994 130 64046
rect 286 63994 329 64046
rect 71 63934 329 63994
rect 71 63882 130 63934
rect 286 63882 329 63934
rect 71 63822 329 63882
rect 71 63770 130 63822
rect 286 63770 329 63822
rect 71 63710 329 63770
rect 71 63658 130 63710
rect 286 63658 329 63710
rect 71 63618 329 63658
rect 71 50658 82 63618
rect 318 50658 329 63618
rect 71 50536 329 50658
rect 71 50484 127 50536
rect 179 50484 239 50536
rect 291 50484 329 50536
rect 71 50424 329 50484
rect 71 50372 127 50424
rect 179 50372 239 50424
rect 291 50372 329 50424
rect 71 50312 329 50372
rect 71 50260 127 50312
rect 179 50260 239 50312
rect 291 50260 329 50312
rect 71 50200 329 50260
rect 71 50148 127 50200
rect 179 50148 239 50200
rect 291 50148 329 50200
rect 71 50088 329 50148
rect 71 50036 127 50088
rect 179 50036 239 50088
rect 291 50036 329 50088
rect 71 49976 329 50036
rect 71 49924 127 49976
rect 179 49924 239 49976
rect 291 49924 329 49976
rect 71 49864 329 49924
rect 71 49812 127 49864
rect 179 49812 239 49864
rect 291 49812 329 49864
rect 71 49752 329 49812
rect 71 49700 127 49752
rect 179 49700 239 49752
rect 291 49700 329 49752
rect 71 49640 329 49700
rect 71 49588 127 49640
rect 179 49588 239 49640
rect 291 49588 329 49640
rect 71 49528 329 49588
rect 71 49476 127 49528
rect 179 49476 239 49528
rect 291 49476 329 49528
rect 71 49416 329 49476
rect 71 49364 127 49416
rect 179 49364 239 49416
rect 291 49364 329 49416
rect 71 49304 329 49364
rect 71 49252 127 49304
rect 179 49252 239 49304
rect 291 49252 329 49304
rect 71 49150 329 49252
rect 71 13276 82 49150
rect 318 13276 329 49150
rect 71 13265 329 13276
rect 375 13151 432 69897
rect -32 13119 127 13151
rect 273 13119 432 13151
rect -32 13108 432 13119
<< via1 >>
rect 130 64890 286 64942
rect 130 64778 286 64830
rect 130 64666 286 64718
rect 130 64554 286 64606
rect 130 64442 286 64494
rect 130 64330 286 64382
rect 130 64218 286 64270
rect 130 64106 286 64158
rect 130 63994 286 64046
rect 130 63882 286 63934
rect 130 63770 286 63822
rect 130 63658 286 63710
rect 127 50484 179 50536
rect 239 50484 291 50536
rect 127 50372 179 50424
rect 239 50372 291 50424
rect 127 50260 179 50312
rect 239 50260 291 50312
rect 127 50148 179 50200
rect 239 50148 291 50200
rect 127 50036 179 50088
rect 239 50036 291 50088
rect 127 49924 179 49976
rect 239 49924 291 49976
rect 127 49812 179 49864
rect 239 49812 291 49864
rect 127 49700 179 49752
rect 239 49700 291 49752
rect 127 49588 179 49640
rect 239 49588 291 49640
rect 127 49476 179 49528
rect 239 49476 291 49528
rect 127 49364 179 49416
rect 239 49364 291 49416
rect 127 49252 179 49304
rect 239 49252 291 49304
<< metal2 >>
rect 118 65000 298 69769
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 118 50600 298 63600
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
rect 118 13275 298 49200
<< via2 >>
rect 128 64942 288 64944
rect 128 64890 130 64942
rect 130 64890 286 64942
rect 286 64890 288 64942
rect 128 64888 288 64890
rect 128 64830 288 64832
rect 128 64778 130 64830
rect 130 64778 286 64830
rect 286 64778 288 64830
rect 128 64776 288 64778
rect 128 64718 288 64720
rect 128 64666 130 64718
rect 130 64666 286 64718
rect 286 64666 288 64718
rect 128 64664 288 64666
rect 128 64606 288 64608
rect 128 64554 130 64606
rect 130 64554 286 64606
rect 286 64554 288 64606
rect 128 64552 288 64554
rect 128 64494 288 64496
rect 128 64442 130 64494
rect 130 64442 286 64494
rect 286 64442 288 64494
rect 128 64440 288 64442
rect 128 64382 288 64384
rect 128 64330 130 64382
rect 130 64330 286 64382
rect 286 64330 288 64382
rect 128 64328 288 64330
rect 128 64270 288 64272
rect 128 64218 130 64270
rect 130 64218 286 64270
rect 286 64218 288 64270
rect 128 64216 288 64218
rect 128 64158 288 64160
rect 128 64106 130 64158
rect 130 64106 286 64158
rect 286 64106 288 64158
rect 128 64104 288 64106
rect 128 64046 288 64048
rect 128 63994 130 64046
rect 130 63994 286 64046
rect 286 63994 288 64046
rect 128 63992 288 63994
rect 128 63934 288 63936
rect 128 63882 130 63934
rect 130 63882 286 63934
rect 286 63882 288 63934
rect 128 63880 288 63882
rect 128 63822 288 63824
rect 128 63770 130 63822
rect 130 63770 286 63822
rect 286 63770 288 63822
rect 128 63768 288 63770
rect 128 63710 288 63712
rect 128 63658 130 63710
rect 130 63658 286 63710
rect 286 63658 288 63710
rect 128 63656 288 63658
rect 125 50536 181 50538
rect 125 50484 127 50536
rect 127 50484 179 50536
rect 179 50484 181 50536
rect 125 50482 181 50484
rect 237 50536 293 50538
rect 237 50484 239 50536
rect 239 50484 291 50536
rect 291 50484 293 50536
rect 237 50482 293 50484
rect 125 50424 181 50426
rect 125 50372 127 50424
rect 127 50372 179 50424
rect 179 50372 181 50424
rect 125 50370 181 50372
rect 237 50424 293 50426
rect 237 50372 239 50424
rect 239 50372 291 50424
rect 291 50372 293 50424
rect 237 50370 293 50372
rect 125 50312 181 50314
rect 125 50260 127 50312
rect 127 50260 179 50312
rect 179 50260 181 50312
rect 125 50258 181 50260
rect 237 50312 293 50314
rect 237 50260 239 50312
rect 239 50260 291 50312
rect 291 50260 293 50312
rect 237 50258 293 50260
rect 125 50200 181 50202
rect 125 50148 127 50200
rect 127 50148 179 50200
rect 179 50148 181 50200
rect 125 50146 181 50148
rect 237 50200 293 50202
rect 237 50148 239 50200
rect 239 50148 291 50200
rect 291 50148 293 50200
rect 237 50146 293 50148
rect 125 50088 181 50090
rect 125 50036 127 50088
rect 127 50036 179 50088
rect 179 50036 181 50088
rect 125 50034 181 50036
rect 237 50088 293 50090
rect 237 50036 239 50088
rect 239 50036 291 50088
rect 291 50036 293 50088
rect 237 50034 293 50036
rect 125 49976 181 49978
rect 125 49924 127 49976
rect 127 49924 179 49976
rect 179 49924 181 49976
rect 125 49922 181 49924
rect 237 49976 293 49978
rect 237 49924 239 49976
rect 239 49924 291 49976
rect 291 49924 293 49976
rect 237 49922 293 49924
rect 125 49864 181 49866
rect 125 49812 127 49864
rect 127 49812 179 49864
rect 179 49812 181 49864
rect 125 49810 181 49812
rect 237 49864 293 49866
rect 237 49812 239 49864
rect 239 49812 291 49864
rect 291 49812 293 49864
rect 237 49810 293 49812
rect 125 49752 181 49754
rect 125 49700 127 49752
rect 127 49700 179 49752
rect 179 49700 181 49752
rect 125 49698 181 49700
rect 237 49752 293 49754
rect 237 49700 239 49752
rect 239 49700 291 49752
rect 291 49700 293 49752
rect 237 49698 293 49700
rect 125 49640 181 49642
rect 125 49588 127 49640
rect 127 49588 179 49640
rect 179 49588 181 49640
rect 125 49586 181 49588
rect 237 49640 293 49642
rect 237 49588 239 49640
rect 239 49588 291 49640
rect 291 49588 293 49640
rect 237 49586 293 49588
rect 125 49528 181 49530
rect 125 49476 127 49528
rect 127 49476 179 49528
rect 179 49476 181 49528
rect 125 49474 181 49476
rect 237 49528 293 49530
rect 237 49476 239 49528
rect 239 49476 291 49528
rect 291 49476 293 49528
rect 237 49474 293 49476
rect 125 49416 181 49418
rect 125 49364 127 49416
rect 127 49364 179 49416
rect 179 49364 181 49416
rect 125 49362 181 49364
rect 237 49416 293 49418
rect 237 49364 239 49416
rect 239 49364 291 49416
rect 291 49364 293 49416
rect 237 49362 293 49364
rect 125 49304 181 49306
rect 125 49252 127 49304
rect 127 49252 179 49304
rect 179 49252 181 49304
rect 125 49250 181 49252
rect 237 49304 293 49306
rect 237 49252 239 49304
rect 239 49252 291 49304
rect 291 49252 293 49304
rect 237 49250 293 49252
<< metal3 >>
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_0
timestamp 1750858719
transform -1 0 48 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_1
timestamp 1750858719
transform 1 0 352 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_40661956134187  M1_PSUB_CDNS_40661956134187_0
timestamp 1750858719
transform 1 0 200 0 -1 13192
box 0 0 1 1
use M1_PSUB_CDNS_40661956134187  M1_PSUB_CDNS_40661956134187_1
timestamp 1750858719
transform 1 0 200 0 1 69873
box 0 0 1 1
use M2_M1_CDNS_40661956134184  M2_M1_CDNS_40661956134184_0
timestamp 1750858719
transform 1 0 208 0 1 64300
box 0 0 1 1
use M2_M1_CDNS_40661956134186  M2_M1_CDNS_40661956134186_0
timestamp 1750858719
transform 1 0 209 0 1 49894
box 0 0 1 1
use M3_M2_CDNS_40661956134183  M3_M2_CDNS_40661956134183_0
timestamp 1750858719
transform 1 0 208 0 1 64300
box 0 0 1 1
use M3_M2_CDNS_40661956134185  M3_M2_CDNS_40661956134185_0
timestamp 1750858719
transform 1 0 209 0 1 49894
box 0 0 1 1
use POLY_FILL  POLY_FILL_0
array 0 0 0 0 351 160
timestamp 1750858719
transform 1 0 82 0 1 13462
box 0 -76 236 84
<< labels >>
rlabel metal3 s 0 63600 400 65000 4 VSS
port 1 nsew ground bidirectional
rlabel metal3 s 0 49200 400 50600 4 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 400 70000
string GDS_END 2921822
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2919750
string LEFclass PAD
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
