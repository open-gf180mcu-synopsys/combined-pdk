magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3440 1660
<< nmos >>
rect 230 210 290 380
rect 340 210 400 380
rect 690 210 750 380
rect 850 210 910 380
rect 1020 210 1080 380
rect 1130 210 1190 380
rect 1300 210 1360 380
rect 1410 210 1470 380
rect 1580 210 1640 380
rect 1690 210 1750 380
rect 1860 210 1920 380
rect 2200 210 2260 380
rect 2550 210 2610 380
rect 2660 210 2720 380
rect 3010 210 3070 380
rect 3180 210 3240 380
<< pmos >>
rect 200 1110 260 1450
rect 370 1110 430 1450
rect 690 1110 750 1450
rect 850 1110 910 1450
rect 1020 1110 1080 1450
rect 1130 1110 1190 1450
rect 1300 1110 1360 1450
rect 1410 1110 1470 1450
rect 1580 1110 1640 1450
rect 1690 1110 1750 1450
rect 1860 1110 1920 1450
rect 2200 1110 2260 1450
rect 2520 1110 2580 1450
rect 2690 1110 2750 1450
rect 3010 1110 3070 1450
rect 3180 1110 3240 1450
<< ndiff >>
rect 120 318 230 380
rect 120 272 152 318
rect 198 272 230 318
rect 120 210 230 272
rect 290 210 340 380
rect 400 318 500 380
rect 400 272 432 318
rect 478 272 500 318
rect 400 210 500 272
rect 590 318 690 380
rect 590 272 612 318
rect 658 272 690 318
rect 590 210 690 272
rect 750 210 850 380
rect 910 318 1020 380
rect 910 272 942 318
rect 988 272 1020 318
rect 910 210 1020 272
rect 1080 210 1130 380
rect 1190 278 1300 380
rect 1190 232 1222 278
rect 1268 232 1300 278
rect 1190 210 1300 232
rect 1360 210 1410 380
rect 1470 318 1580 380
rect 1470 272 1502 318
rect 1548 272 1580 318
rect 1470 210 1580 272
rect 1640 210 1690 380
rect 1750 318 1860 380
rect 1750 272 1782 318
rect 1828 272 1860 318
rect 1750 210 1860 272
rect 1920 318 2020 380
rect 1920 272 1952 318
rect 1998 272 2020 318
rect 1920 210 2020 272
rect 2100 318 2200 380
rect 2100 272 2122 318
rect 2168 272 2200 318
rect 2100 210 2200 272
rect 2260 318 2360 380
rect 2260 272 2292 318
rect 2338 272 2360 318
rect 2260 210 2360 272
rect 2450 318 2550 380
rect 2450 272 2472 318
rect 2518 272 2550 318
rect 2450 210 2550 272
rect 2610 210 2660 380
rect 2720 318 2820 380
rect 2720 272 2752 318
rect 2798 272 2820 318
rect 2720 210 2820 272
rect 2910 318 3010 380
rect 2910 272 2932 318
rect 2978 272 3010 318
rect 2910 210 3010 272
rect 3070 318 3180 380
rect 3070 272 3102 318
rect 3148 272 3180 318
rect 3070 210 3180 272
rect 3240 318 3340 380
rect 3240 272 3272 318
rect 3318 272 3340 318
rect 3240 210 3340 272
<< pdiff >>
rect 90 1425 200 1450
rect 90 1285 122 1425
rect 168 1285 200 1425
rect 90 1110 200 1285
rect 260 1425 370 1450
rect 260 1285 292 1425
rect 338 1285 370 1425
rect 260 1110 370 1285
rect 430 1425 530 1450
rect 430 1285 462 1425
rect 508 1285 530 1425
rect 430 1110 530 1285
rect 590 1397 690 1450
rect 590 1163 612 1397
rect 658 1163 690 1397
rect 590 1110 690 1163
rect 750 1110 850 1450
rect 910 1397 1020 1450
rect 910 1163 942 1397
rect 988 1163 1020 1397
rect 910 1110 1020 1163
rect 1080 1110 1130 1450
rect 1190 1397 1300 1450
rect 1190 1163 1222 1397
rect 1268 1163 1300 1397
rect 1190 1110 1300 1163
rect 1360 1110 1410 1450
rect 1470 1425 1580 1450
rect 1470 1285 1502 1425
rect 1548 1285 1580 1425
rect 1470 1110 1580 1285
rect 1640 1110 1690 1450
rect 1750 1425 1860 1450
rect 1750 1285 1782 1425
rect 1828 1285 1860 1425
rect 1750 1110 1860 1285
rect 1920 1397 2020 1450
rect 1920 1163 1952 1397
rect 1998 1163 2020 1397
rect 1920 1110 2020 1163
rect 2100 1397 2200 1450
rect 2100 1163 2122 1397
rect 2168 1163 2200 1397
rect 2100 1110 2200 1163
rect 2260 1397 2360 1450
rect 2260 1163 2292 1397
rect 2338 1163 2360 1397
rect 2260 1110 2360 1163
rect 2420 1430 2520 1450
rect 2420 1290 2442 1430
rect 2488 1290 2520 1430
rect 2420 1110 2520 1290
rect 2580 1428 2690 1450
rect 2580 1382 2612 1428
rect 2658 1382 2690 1428
rect 2580 1110 2690 1382
rect 2750 1388 2850 1450
rect 2750 1342 2782 1388
rect 2828 1342 2850 1388
rect 2750 1110 2850 1342
rect 2910 1397 3010 1450
rect 2910 1163 2932 1397
rect 2978 1163 3010 1397
rect 2910 1110 3010 1163
rect 3070 1397 3180 1450
rect 3070 1163 3102 1397
rect 3148 1163 3180 1397
rect 3070 1110 3180 1163
rect 3240 1397 3340 1450
rect 3240 1163 3272 1397
rect 3318 1163 3340 1397
rect 3240 1110 3340 1163
<< ndiffc >>
rect 152 272 198 318
rect 432 272 478 318
rect 612 272 658 318
rect 942 272 988 318
rect 1222 232 1268 278
rect 1502 272 1548 318
rect 1782 272 1828 318
rect 1952 272 1998 318
rect 2122 272 2168 318
rect 2292 272 2338 318
rect 2472 272 2518 318
rect 2752 272 2798 318
rect 2932 272 2978 318
rect 3102 272 3148 318
rect 3272 272 3318 318
<< pdiffc >>
rect 122 1285 168 1425
rect 292 1285 338 1425
rect 462 1285 508 1425
rect 612 1163 658 1397
rect 942 1163 988 1397
rect 1222 1163 1268 1397
rect 1502 1285 1548 1425
rect 1782 1285 1828 1425
rect 1952 1163 1998 1397
rect 2122 1163 2168 1397
rect 2292 1163 2338 1397
rect 2442 1290 2488 1430
rect 2612 1382 2658 1428
rect 2782 1342 2828 1388
rect 2932 1163 2978 1397
rect 3102 1163 3148 1397
rect 3272 1163 3318 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
rect 980 118 1130 140
rect 980 72 1032 118
rect 1078 72 1130 118
rect 980 50 1130 72
rect 1210 118 1360 140
rect 1210 72 1262 118
rect 1308 72 1360 118
rect 1210 50 1360 72
rect 1440 118 1590 140
rect 1440 72 1492 118
rect 1538 72 1590 118
rect 1440 50 1590 72
rect 1670 118 1820 140
rect 1670 72 1722 118
rect 1768 72 1820 118
rect 1670 50 1820 72
rect 1900 118 2050 140
rect 1900 72 1952 118
rect 1998 72 2050 118
rect 1900 50 2050 72
rect 2130 118 2280 140
rect 2130 72 2182 118
rect 2228 72 2280 118
rect 2130 50 2280 72
rect 2360 118 2510 140
rect 2360 72 2412 118
rect 2458 72 2510 118
rect 2360 50 2510 72
rect 2590 118 2740 140
rect 2590 72 2642 118
rect 2688 72 2740 118
rect 2590 50 2740 72
rect 2820 118 2970 140
rect 2820 72 2872 118
rect 2918 72 2970 118
rect 2820 50 2970 72
rect 3050 118 3200 140
rect 3050 72 3102 118
rect 3148 72 3200 118
rect 3050 50 3200 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
rect 980 1588 1130 1610
rect 980 1542 1032 1588
rect 1078 1542 1130 1588
rect 980 1520 1130 1542
rect 1210 1588 1360 1610
rect 1210 1542 1262 1588
rect 1308 1542 1360 1588
rect 1210 1520 1360 1542
rect 1440 1588 1590 1610
rect 1440 1542 1492 1588
rect 1538 1542 1590 1588
rect 1440 1520 1590 1542
rect 1670 1588 1820 1610
rect 1670 1542 1722 1588
rect 1768 1542 1820 1588
rect 1670 1520 1820 1542
rect 1900 1588 2050 1610
rect 1900 1542 1952 1588
rect 1998 1542 2050 1588
rect 1900 1520 2050 1542
rect 2130 1588 2280 1610
rect 2130 1542 2182 1588
rect 2228 1542 2280 1588
rect 2130 1520 2280 1542
rect 2360 1588 2510 1610
rect 2360 1542 2412 1588
rect 2458 1542 2510 1588
rect 2360 1520 2510 1542
rect 2590 1588 2740 1610
rect 2590 1542 2642 1588
rect 2688 1542 2740 1588
rect 2590 1520 2740 1542
rect 2820 1588 2970 1610
rect 2820 1542 2872 1588
rect 2918 1542 2970 1588
rect 2820 1520 2970 1542
rect 3050 1588 3200 1610
rect 3050 1542 3102 1588
rect 3148 1542 3200 1588
rect 3050 1520 3200 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
rect 1032 72 1078 118
rect 1262 72 1308 118
rect 1492 72 1538 118
rect 1722 72 1768 118
rect 1952 72 1998 118
rect 2182 72 2228 118
rect 2412 72 2458 118
rect 2642 72 2688 118
rect 2872 72 2918 118
rect 3102 72 3148 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
rect 1032 1542 1078 1588
rect 1262 1542 1308 1588
rect 1492 1542 1538 1588
rect 1722 1542 1768 1588
rect 1952 1542 1998 1588
rect 2182 1542 2228 1588
rect 2412 1542 2458 1588
rect 2642 1542 2688 1588
rect 2872 1542 2918 1588
rect 3102 1542 3148 1588
<< polysilicon >>
rect 200 1450 260 1500
rect 370 1450 430 1500
rect 690 1450 750 1500
rect 850 1450 910 1500
rect 1020 1450 1080 1500
rect 1130 1450 1190 1500
rect 1300 1450 1360 1500
rect 1410 1450 1470 1500
rect 1580 1450 1640 1500
rect 1690 1450 1750 1500
rect 1860 1450 1920 1500
rect 2200 1450 2260 1500
rect 2520 1450 2580 1500
rect 2690 1450 2750 1500
rect 3010 1450 3070 1500
rect 3180 1450 3240 1500
rect 200 930 260 1110
rect 200 903 320 930
rect 200 857 227 903
rect 273 857 320 903
rect 200 830 320 857
rect 200 470 260 830
rect 370 800 430 1110
rect 690 800 750 1110
rect 850 930 910 1110
rect 850 903 950 930
rect 850 857 877 903
rect 923 857 950 903
rect 850 830 950 857
rect 370 773 510 800
rect 370 727 427 773
rect 473 727 510 773
rect 370 700 510 727
rect 690 773 810 800
rect 690 727 737 773
rect 783 727 810 773
rect 690 700 810 727
rect 370 470 430 700
rect 200 430 290 470
rect 230 380 290 430
rect 340 430 430 470
rect 340 380 400 430
rect 690 380 750 700
rect 1020 660 1080 1110
rect 1130 1060 1190 1110
rect 1300 1060 1360 1110
rect 1130 1033 1360 1060
rect 1130 990 1167 1033
rect 1140 987 1167 990
rect 1213 990 1360 1033
rect 1213 987 1240 990
rect 1140 940 1240 987
rect 1410 660 1470 1110
rect 1580 930 1640 1110
rect 1540 903 1640 930
rect 1540 857 1567 903
rect 1613 857 1640 903
rect 1540 830 1640 857
rect 1690 800 1750 1110
rect 1860 930 1920 1110
rect 1860 903 1960 930
rect 1860 857 1887 903
rect 1933 857 1960 903
rect 1860 830 1960 857
rect 1680 773 1780 800
rect 1680 727 1707 773
rect 1753 727 1780 773
rect 1680 700 1780 727
rect 1540 660 1640 670
rect 850 643 1640 660
rect 850 600 1567 643
rect 850 380 910 600
rect 1540 597 1567 600
rect 1613 597 1640 643
rect 1540 570 1640 597
rect 980 513 1080 540
rect 1140 520 1240 540
rect 980 467 1007 513
rect 1053 467 1080 513
rect 980 440 1080 467
rect 1020 380 1080 440
rect 1130 513 1360 520
rect 1130 467 1167 513
rect 1213 467 1360 513
rect 1130 440 1360 467
rect 1130 380 1190 440
rect 1300 380 1360 440
rect 1410 503 1510 530
rect 1410 457 1437 503
rect 1483 457 1510 503
rect 1410 430 1510 457
rect 1410 380 1470 430
rect 1580 380 1640 570
rect 1690 380 1750 700
rect 1860 380 1920 830
rect 2200 670 2260 1110
rect 2200 643 2340 670
rect 2200 597 2267 643
rect 2313 597 2340 643
rect 2200 570 2340 597
rect 2200 380 2260 570
rect 2520 530 2580 1110
rect 2690 930 2750 1110
rect 2630 903 2750 930
rect 2630 857 2677 903
rect 2723 857 2750 903
rect 2630 830 2750 857
rect 2440 503 2580 530
rect 2440 457 2477 503
rect 2523 470 2580 503
rect 2690 470 2750 830
rect 3010 670 3070 1110
rect 3180 930 3240 1110
rect 3120 903 3240 930
rect 3120 857 3147 903
rect 3193 857 3240 903
rect 3120 830 3240 857
rect 2950 643 3070 670
rect 2950 597 2997 643
rect 3043 597 3070 643
rect 2950 570 3070 597
rect 2523 457 2610 470
rect 2440 430 2610 457
rect 2550 380 2610 430
rect 2660 430 2750 470
rect 2660 380 2720 430
rect 3010 380 3070 570
rect 3180 380 3240 830
rect 230 160 290 210
rect 340 160 400 210
rect 690 160 750 210
rect 850 160 910 210
rect 1020 160 1080 210
rect 1130 160 1190 210
rect 1300 160 1360 210
rect 1410 160 1470 210
rect 1580 160 1640 210
rect 1690 160 1750 210
rect 1860 160 1920 210
rect 2200 160 2260 210
rect 2550 160 2610 210
rect 2660 160 2720 210
rect 3010 160 3070 210
rect 3180 160 3240 210
<< polycontact >>
rect 227 857 273 903
rect 877 857 923 903
rect 427 727 473 773
rect 737 727 783 773
rect 1167 987 1213 1033
rect 1567 857 1613 903
rect 1887 857 1933 903
rect 1707 727 1753 773
rect 1567 597 1613 643
rect 1007 467 1053 513
rect 1167 467 1213 513
rect 1437 457 1483 503
rect 2267 597 2313 643
rect 2677 857 2723 903
rect 2477 457 2523 503
rect 3147 857 3193 903
rect 2997 597 3043 643
<< metal1 >>
rect 0 1588 3440 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1032 1588
rect 1078 1542 1262 1588
rect 1308 1542 1492 1588
rect 1538 1542 1722 1588
rect 1768 1542 1952 1588
rect 1998 1542 2182 1588
rect 2228 1542 2412 1588
rect 2458 1542 2642 1588
rect 2688 1542 2872 1588
rect 2918 1542 3102 1588
rect 3148 1542 3440 1588
rect 0 1520 3440 1542
rect 120 1425 170 1450
rect 120 1285 122 1425
rect 168 1285 170 1425
rect 120 1210 170 1285
rect 290 1425 340 1520
rect 290 1285 292 1425
rect 338 1285 340 1425
rect 290 1260 340 1285
rect 460 1425 510 1450
rect 460 1285 462 1425
rect 508 1285 510 1425
rect 460 1210 510 1285
rect 120 1160 510 1210
rect 610 1397 660 1520
rect 610 1163 612 1397
rect 658 1163 660 1397
rect 150 910 200 1160
rect 610 1110 660 1163
rect 940 1397 990 1450
rect 940 1163 942 1397
rect 988 1163 990 1397
rect 940 1060 990 1163
rect 1220 1397 1270 1520
rect 1220 1163 1222 1397
rect 1268 1163 1270 1397
rect 1500 1425 1550 1450
rect 1500 1285 1502 1425
rect 1548 1285 1550 1425
rect 1500 1260 1550 1285
rect 1780 1425 1830 1520
rect 1780 1285 1782 1425
rect 1828 1285 1830 1425
rect 1780 1260 1830 1285
rect 1950 1397 2000 1450
rect 1220 1110 1270 1163
rect 1320 1210 1550 1260
rect 610 1010 990 1060
rect 1140 1033 1240 1040
rect 150 906 300 910
rect 150 854 224 906
rect 276 854 300 906
rect 150 850 300 854
rect 150 520 200 850
rect 610 780 660 1010
rect 1140 987 1167 1033
rect 1213 987 1240 1033
rect 1140 980 1240 987
rect 850 906 1080 910
rect 850 903 1004 906
rect 850 857 877 903
rect 923 857 1004 903
rect 850 854 1004 857
rect 1056 854 1080 906
rect 850 850 1080 854
rect 400 776 660 780
rect 400 724 424 776
rect 476 724 660 776
rect 400 720 660 724
rect 710 776 810 780
rect 710 724 734 776
rect 786 724 810 776
rect 710 720 810 724
rect 420 520 470 530
rect 610 520 660 720
rect 1000 520 1060 850
rect 1160 520 1220 980
rect 1320 760 1370 1210
rect 1950 1163 1952 1397
rect 1998 1163 2000 1397
rect 1670 1036 1770 1040
rect 1670 984 1694 1036
rect 1746 984 1770 1036
rect 1670 980 1770 984
rect 1950 1020 2000 1163
rect 2120 1397 2170 1450
rect 2120 1163 2122 1397
rect 2168 1163 2170 1397
rect 2120 1140 2170 1163
rect 1310 710 1370 760
rect 1430 906 1640 910
rect 1430 854 1564 906
rect 1616 854 1640 906
rect 1430 850 1640 854
rect 150 516 500 520
rect 150 464 424 516
rect 476 464 500 516
rect 610 470 810 520
rect 150 460 500 464
rect 150 318 200 460
rect 420 450 470 460
rect 730 380 810 470
rect 980 513 1080 520
rect 980 467 1007 513
rect 1053 467 1080 513
rect 980 460 1080 467
rect 1140 516 1240 520
rect 1140 464 1164 516
rect 1216 464 1240 516
rect 1140 460 1240 464
rect 1310 390 1360 710
rect 1430 510 1490 850
rect 1690 780 1750 980
rect 1950 970 2060 1020
rect 1860 906 1960 910
rect 1860 854 1884 906
rect 1936 854 1960 906
rect 1860 850 1960 854
rect 2010 780 2060 970
rect 1680 776 1780 780
rect 1680 724 1704 776
rect 1756 724 1780 776
rect 1680 720 1780 724
rect 1950 730 2060 780
rect 2110 910 2170 1140
rect 2290 1397 2340 1520
rect 2290 1163 2292 1397
rect 2338 1163 2340 1397
rect 2440 1430 2490 1450
rect 2440 1290 2442 1430
rect 2488 1310 2490 1430
rect 2610 1428 2660 1520
rect 2610 1382 2612 1428
rect 2658 1382 2660 1428
rect 2610 1360 2660 1382
rect 2780 1388 2830 1450
rect 2780 1342 2782 1388
rect 2828 1342 2830 1388
rect 2780 1310 2830 1342
rect 2488 1290 2830 1310
rect 2440 1260 2830 1290
rect 2930 1397 2980 1450
rect 2290 1110 2340 1163
rect 2930 1163 2932 1397
rect 2978 1163 2980 1397
rect 2470 1040 2530 1060
rect 2810 1040 2870 1060
rect 2470 1036 2870 1040
rect 2470 984 2474 1036
rect 2526 984 2814 1036
rect 2866 984 2870 1036
rect 2470 980 2870 984
rect 2470 960 2530 980
rect 2110 906 2180 910
rect 2110 854 2114 906
rect 2166 854 2180 906
rect 2110 850 2180 854
rect 2650 906 2750 910
rect 2650 854 2674 906
rect 2726 854 2750 906
rect 2650 850 2750 854
rect 1540 646 1640 650
rect 1540 594 1564 646
rect 1616 594 1640 646
rect 1540 590 1640 594
rect 1950 646 2010 730
rect 1950 594 1954 646
rect 2006 594 2010 646
rect 1950 570 2010 594
rect 1410 503 1510 510
rect 1410 457 1437 503
rect 1483 457 1510 503
rect 1410 450 1510 457
rect 1310 386 1580 390
rect 150 272 152 318
rect 198 272 200 318
rect 150 210 200 272
rect 430 318 480 380
rect 430 272 432 318
rect 478 272 480 318
rect 430 140 480 272
rect 610 318 660 380
rect 730 330 990 380
rect 1310 340 1504 386
rect 610 272 612 318
rect 658 272 660 318
rect 610 140 660 272
rect 940 318 990 330
rect 940 272 942 318
rect 988 272 990 318
rect 1500 334 1504 340
rect 1556 334 1580 386
rect 1500 330 1580 334
rect 1500 318 1550 330
rect 940 210 990 272
rect 1220 278 1270 300
rect 1220 232 1222 278
rect 1268 232 1270 278
rect 1220 140 1270 232
rect 1500 272 1502 318
rect 1548 272 1550 318
rect 1500 210 1550 272
rect 1780 318 1830 380
rect 1780 272 1782 318
rect 1828 272 1830 318
rect 1780 140 1830 272
rect 1950 318 2000 570
rect 2110 360 2170 850
rect 2810 650 2870 980
rect 2930 910 2980 1163
rect 3100 1397 3150 1520
rect 3100 1163 3102 1397
rect 3148 1163 3150 1397
rect 3100 1110 3150 1163
rect 3270 1397 3320 1450
rect 3270 1163 3272 1397
rect 3318 1163 3320 1397
rect 3270 1050 3320 1163
rect 3270 1036 3370 1050
rect 3270 984 3294 1036
rect 3346 984 3370 1036
rect 3270 980 3370 984
rect 3270 970 3360 980
rect 2930 906 3220 910
rect 2930 854 3144 906
rect 3196 854 3220 906
rect 2930 850 3220 854
rect 2240 646 2340 650
rect 2240 594 2264 646
rect 2316 594 2340 646
rect 2240 590 2340 594
rect 2750 646 3070 650
rect 2750 594 2994 646
rect 3046 594 3070 646
rect 2750 590 3070 594
rect 2450 506 2550 510
rect 2450 454 2474 506
rect 2526 454 2550 506
rect 2450 450 2550 454
rect 1950 272 1952 318
rect 1998 272 2000 318
rect 1950 210 2000 272
rect 2120 318 2170 360
rect 2120 272 2122 318
rect 2168 272 2170 318
rect 2120 210 2170 272
rect 2290 318 2340 380
rect 2290 272 2292 318
rect 2338 272 2340 318
rect 2290 140 2340 272
rect 2470 318 2520 380
rect 2470 272 2472 318
rect 2518 272 2520 318
rect 2470 140 2520 272
rect 2750 318 2800 590
rect 3150 480 3200 850
rect 2750 272 2752 318
rect 2798 272 2800 318
rect 2750 210 2800 272
rect 2930 430 3200 480
rect 2930 318 2980 430
rect 2930 272 2932 318
rect 2978 272 2980 318
rect 2930 210 2980 272
rect 3100 318 3150 380
rect 3100 272 3102 318
rect 3148 272 3150 318
rect 3100 140 3150 272
rect 3270 318 3320 970
rect 3270 272 3272 318
rect 3318 272 3320 318
rect 3270 210 3320 272
rect 0 118 3440 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1032 118
rect 1078 72 1262 118
rect 1308 72 1492 118
rect 1538 72 1722 118
rect 1768 72 1952 118
rect 1998 72 2182 118
rect 2228 72 2412 118
rect 2458 72 2642 118
rect 2688 72 2872 118
rect 2918 72 3102 118
rect 3148 72 3440 118
rect 0 0 3440 72
<< via1 >>
rect 224 903 276 906
rect 224 857 227 903
rect 227 857 273 903
rect 273 857 276 903
rect 224 854 276 857
rect 1004 854 1056 906
rect 424 773 476 776
rect 424 727 427 773
rect 427 727 473 773
rect 473 727 476 773
rect 424 724 476 727
rect 734 773 786 776
rect 734 727 737 773
rect 737 727 783 773
rect 783 727 786 773
rect 734 724 786 727
rect 1694 984 1746 1036
rect 1564 903 1616 906
rect 1564 857 1567 903
rect 1567 857 1613 903
rect 1613 857 1616 903
rect 1564 854 1616 857
rect 424 464 476 516
rect 1164 513 1216 516
rect 1164 467 1167 513
rect 1167 467 1213 513
rect 1213 467 1216 513
rect 1164 464 1216 467
rect 1884 903 1936 906
rect 1884 857 1887 903
rect 1887 857 1933 903
rect 1933 857 1936 903
rect 1884 854 1936 857
rect 1704 773 1756 776
rect 1704 727 1707 773
rect 1707 727 1753 773
rect 1753 727 1756 773
rect 1704 724 1756 727
rect 2474 984 2526 1036
rect 2814 984 2866 1036
rect 2114 854 2166 906
rect 2674 903 2726 906
rect 2674 857 2677 903
rect 2677 857 2723 903
rect 2723 857 2726 903
rect 2674 854 2726 857
rect 1564 643 1616 646
rect 1564 597 1567 643
rect 1567 597 1613 643
rect 1613 597 1616 643
rect 1564 594 1616 597
rect 1954 594 2006 646
rect 1504 334 1556 386
rect 3294 984 3346 1036
rect 3144 903 3196 906
rect 3144 857 3147 903
rect 3147 857 3193 903
rect 3193 857 3196 903
rect 3144 854 3196 857
rect 2264 643 2316 646
rect 2264 597 2267 643
rect 2267 597 2313 643
rect 2313 597 2316 643
rect 2264 594 2316 597
rect 2994 643 3046 646
rect 2994 597 2997 643
rect 2997 597 3043 643
rect 3043 597 3046 643
rect 2994 594 3046 597
rect 2474 503 2526 506
rect 2474 457 2477 503
rect 2477 457 2523 503
rect 2523 457 2526 503
rect 2474 454 2526 457
<< metal2 >>
rect 220 1110 2730 1170
rect 220 920 280 1110
rect 1680 1040 1760 1050
rect 2460 1040 2540 1050
rect 1670 1036 2550 1040
rect 1670 984 1694 1036
rect 1746 984 2474 1036
rect 2526 984 2550 1036
rect 1670 980 2550 984
rect 1680 970 1760 980
rect 2460 970 2540 980
rect 2670 920 2730 1110
rect 2790 1036 2890 1050
rect 3280 1040 3360 1050
rect 2790 984 2814 1036
rect 2866 984 2890 1036
rect 2790 970 2890 984
rect 3270 1036 3370 1040
rect 3270 984 3294 1036
rect 3346 984 3370 1036
rect 3270 980 3370 984
rect 3280 970 3360 980
rect 200 906 300 920
rect 200 854 224 906
rect 276 854 300 906
rect 200 840 300 854
rect 980 910 1070 920
rect 1540 910 1640 920
rect 1870 910 1950 920
rect 2100 910 2180 920
rect 980 906 2190 910
rect 980 854 1004 906
rect 1056 854 1564 906
rect 1616 854 1884 906
rect 1936 854 2114 906
rect 2166 854 2190 906
rect 980 850 2190 854
rect 2650 906 2750 920
rect 3130 910 3210 920
rect 2650 854 2674 906
rect 2726 854 2750 906
rect 980 840 1070 850
rect 1540 840 1640 850
rect 1870 840 1950 850
rect 2100 840 2180 850
rect 2650 840 2750 854
rect 3120 906 3220 910
rect 3120 854 3144 906
rect 3196 854 3220 906
rect 3120 850 3220 854
rect 3130 840 3210 850
rect 400 776 500 790
rect 400 724 424 776
rect 476 724 500 776
rect 400 710 500 724
rect 710 776 810 790
rect 1690 780 1770 790
rect 710 724 734 776
rect 786 724 810 776
rect 710 710 810 724
rect 1680 776 1780 780
rect 1680 724 1704 776
rect 1756 724 1780 776
rect 1680 720 1780 724
rect 1690 710 1770 720
rect 1550 650 1630 660
rect 1940 650 2020 660
rect 2250 650 2330 660
rect 2980 650 3060 660
rect 1540 646 2040 650
rect 1540 594 1564 646
rect 1616 594 1954 646
rect 2006 594 2040 646
rect 1540 590 2040 594
rect 2240 646 2340 650
rect 2240 594 2264 646
rect 2316 594 2340 646
rect 2240 590 2340 594
rect 2910 646 3070 650
rect 2910 594 2994 646
rect 3046 594 3070 646
rect 2910 590 3070 594
rect 1550 580 1630 590
rect 1940 580 2020 590
rect 2250 580 2330 590
rect 2980 580 3060 590
rect 400 520 500 530
rect 1150 520 1230 530
rect 400 516 1240 520
rect 400 464 424 516
rect 476 464 1164 516
rect 1216 464 1240 516
rect 400 460 1240 464
rect 2450 506 2550 520
rect 400 450 500 460
rect 1150 450 1230 460
rect 2450 454 2474 506
rect 2526 454 2550 506
rect 2450 440 2550 454
rect 1490 390 1570 400
rect 2450 390 2530 440
rect 1480 386 2530 390
rect 1480 334 1504 386
rect 1556 334 2530 386
rect 1480 330 2530 334
rect 1490 320 1570 330
<< labels >>
rlabel via1 s 734 724 786 776 4 D
port 1 nsew signal input
rlabel via1 s 3294 984 3346 1036 4 Q
port 2 nsew signal output
rlabel via1 s 3144 854 3196 906 4 QN
port 3 nsew signal output
rlabel via1 s 2264 594 2316 646 4 CLK
port 4 nsew clock input
rlabel via1 s 2674 854 2726 906 4 SN
port 5 nsew signal output
rlabel metal1 s 290 1260 340 1660 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 430 0 480 380 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 610 1110 660 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1220 1110 1270 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1780 1260 1830 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2290 1110 2340 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2610 1360 2660 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3100 1110 3150 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3440 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 0 660 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1220 0 1270 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1780 0 1830 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2290 0 2340 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2470 0 2520 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3100 0 3150 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3440 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal2 s 2250 580 2330 660 1 CLK
port 4 nsew clock input
rlabel metal2 s 2240 590 2340 650 1 CLK
port 4 nsew clock input
rlabel metal1 s 2240 590 2340 650 1 CLK
port 4 nsew clock input
rlabel metal2 s 710 710 810 790 1 D
port 1 nsew signal input
rlabel metal1 s 710 720 810 780 1 D
port 1 nsew signal input
rlabel metal2 s 3280 970 3360 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3270 980 3370 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 3270 210 3320 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 3270 970 3360 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 3270 980 3370 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3130 840 3210 920 1 QN
port 3 nsew signal output
rlabel metal2 s 3120 850 3220 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2930 210 2980 480 1 QN
port 3 nsew signal output
rlabel metal1 s 2930 850 2980 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 2930 430 3200 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3150 430 3200 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2930 850 3220 910 1 QN
port 3 nsew signal output
rlabel via1 s 1164 464 1216 516 1 SN
port 5 nsew signal output
rlabel via1 s 424 464 476 516 1 SN
port 5 nsew signal output
rlabel via1 s 224 854 276 906 1 SN
port 5 nsew signal output
rlabel metal2 s 400 450 500 530 1 SN
port 5 nsew signal output
rlabel metal2 s 1150 450 1230 530 1 SN
port 5 nsew signal output
rlabel metal2 s 400 460 1240 520 1 SN
port 5 nsew signal output
rlabel metal2 s 220 840 280 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 200 840 300 920 1 SN
port 5 nsew signal output
rlabel metal2 s 2670 840 2730 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 220 1110 2730 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 2650 840 2750 920 1 SN
port 5 nsew signal output
rlabel metal1 s 120 1160 170 1450 1 SN
port 5 nsew signal output
rlabel metal1 s 150 210 200 1210 1 SN
port 5 nsew signal output
rlabel metal1 s 150 850 300 910 1 SN
port 5 nsew signal output
rlabel metal1 s 120 1160 510 1210 1 SN
port 5 nsew signal output
rlabel metal1 s 420 450 470 530 1 SN
port 5 nsew signal output
rlabel metal1 s 150 460 500 520 1 SN
port 5 nsew signal output
rlabel metal1 s 460 1160 510 1450 1 SN
port 5 nsew signal output
rlabel metal1 s 1160 460 1220 1040 1 SN
port 5 nsew signal output
rlabel metal1 s 1140 460 1240 520 1 SN
port 5 nsew signal output
rlabel metal1 s 1140 980 1240 1040 1 SN
port 5 nsew signal output
rlabel metal1 s 2650 850 2750 910 1 SN
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3440 1660
string GDS_END 315392
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 290028
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
