magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 7254 870
<< pwell >>
rect -86 -86 7254 352
<< metal1 >>
rect 0 724 7168 844
rect 353 498 399 724
rect 49 60 95 211
rect 801 498 847 724
rect 497 60 543 211
rect 1249 498 1295 724
rect 945 60 991 211
rect 1697 498 1743 724
rect 1393 60 1439 211
rect 2145 498 2191 724
rect 1841 60 1887 211
rect 2593 498 2639 724
rect 2289 60 2335 211
rect 3041 498 3087 724
rect 2737 60 2783 211
rect 3489 498 3535 724
rect 3185 60 3231 211
rect 3937 498 3983 724
rect 3633 60 3679 211
rect 4385 498 4431 724
rect 4081 60 4127 211
rect 4833 498 4879 724
rect 4529 60 4575 211
rect 5281 498 5327 724
rect 4977 60 5023 211
rect 5729 498 5775 724
rect 5425 60 5471 211
rect 6177 498 6223 724
rect 5873 60 5919 211
rect 6625 498 6671 724
rect 6321 60 6367 211
rect 7073 498 7119 724
rect 6769 60 6815 211
rect 0 -60 7168 60
<< obsm1 >>
rect 49 311 95 678
rect 146 392 399 438
rect 49 265 304 311
rect 353 106 399 392
rect 497 311 543 678
rect 594 392 847 438
rect 497 265 752 311
rect 801 106 847 392
rect 945 311 991 678
rect 1042 392 1295 438
rect 945 265 1200 311
rect 1249 106 1295 392
rect 1393 311 1439 678
rect 1490 392 1743 438
rect 1393 265 1648 311
rect 1697 106 1743 392
rect 1841 311 1887 678
rect 1938 392 2191 438
rect 1841 265 2096 311
rect 2145 106 2191 392
rect 2289 311 2335 678
rect 2386 392 2639 438
rect 2289 265 2544 311
rect 2593 106 2639 392
rect 2737 311 2783 678
rect 2834 392 3087 438
rect 2737 265 2992 311
rect 3041 106 3087 392
rect 3185 311 3231 678
rect 3282 392 3535 438
rect 3185 265 3440 311
rect 3489 106 3535 392
rect 3633 311 3679 678
rect 3730 392 3983 438
rect 3633 265 3888 311
rect 3937 106 3983 392
rect 4081 311 4127 678
rect 4178 392 4431 438
rect 4081 265 4336 311
rect 4385 106 4431 392
rect 4529 311 4575 678
rect 4626 392 4879 438
rect 4529 265 4784 311
rect 4833 106 4879 392
rect 4977 311 5023 678
rect 5074 392 5327 438
rect 4977 265 5232 311
rect 5281 106 5327 392
rect 5425 311 5471 678
rect 5522 392 5775 438
rect 5425 265 5680 311
rect 5729 106 5775 392
rect 5873 311 5919 678
rect 5970 392 6223 438
rect 5873 265 6128 311
rect 6177 106 6223 392
rect 6321 311 6367 678
rect 6418 392 6671 438
rect 6321 265 6576 311
rect 6625 106 6671 392
rect 6769 311 6815 678
rect 6866 392 7119 438
rect 6769 265 7024 311
rect 7073 106 7119 392
<< labels >>
rlabel metal1 s 7073 498 7119 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6625 498 6671 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 6177 498 6223 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5729 498 5775 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 5281 498 5327 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4833 498 4879 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 4385 498 4431 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3937 498 3983 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3489 498 3535 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3041 498 3087 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2593 498 2639 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2145 498 2191 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 498 1743 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 498 1295 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 498 847 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 724 7168 844 6 VDD
port 1 nsew power bidirectional abutment
rlabel nwell s -86 352 7254 870 6 VNW
port 2 nsew power bidirectional
rlabel pwell s -86 -86 7254 352 6 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 0 -60 7168 60 8 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6769 60 6815 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6321 60 6367 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5873 60 5919 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5425 60 5471 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4977 60 5023 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 60 4575 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4081 60 4127 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3633 60 3679 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3185 60 3231 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2737 60 2783 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 211 6 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 7168 784
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 421994
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 402914
<< end >>
