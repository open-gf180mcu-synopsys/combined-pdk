magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3740 1660
<< nmos >>
rect 190 210 250 380
rect 540 210 600 380
rect 710 210 770 380
rect 820 210 880 380
rect 1170 210 1230 380
rect 1330 210 1390 380
rect 1500 210 1560 380
rect 1610 210 1670 380
rect 1780 210 1840 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2170 210 2230 380
rect 2340 210 2400 380
rect 2690 210 2750 380
rect 2800 210 2860 380
rect 2970 210 3030 380
rect 3320 210 3380 380
rect 3490 210 3550 380
<< pmos >>
rect 190 1110 250 1450
rect 510 1110 570 1450
rect 680 1110 740 1450
rect 850 1110 910 1450
rect 1170 1110 1230 1450
rect 1330 1110 1390 1450
rect 1500 1110 1560 1450
rect 1610 1110 1670 1450
rect 1780 1110 1840 1450
rect 1890 1110 1950 1450
rect 2060 1110 2120 1450
rect 2170 1110 2230 1450
rect 2340 1110 2400 1450
rect 2660 1110 2720 1450
rect 2830 1110 2890 1450
rect 3000 1110 3060 1450
rect 3320 1110 3380 1450
rect 3490 1110 3550 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 440 318 540 380
rect 440 272 462 318
rect 508 272 540 318
rect 440 210 540 272
rect 600 318 710 380
rect 600 272 632 318
rect 678 272 710 318
rect 600 210 710 272
rect 770 210 820 380
rect 880 318 980 380
rect 880 272 912 318
rect 958 272 980 318
rect 880 210 980 272
rect 1070 318 1170 380
rect 1070 272 1092 318
rect 1138 272 1170 318
rect 1070 210 1170 272
rect 1230 210 1330 380
rect 1390 318 1500 380
rect 1390 272 1422 318
rect 1468 272 1500 318
rect 1390 210 1500 272
rect 1560 210 1610 380
rect 1670 278 1780 380
rect 1670 232 1702 278
rect 1748 232 1780 278
rect 1670 210 1780 232
rect 1840 210 1890 380
rect 1950 318 2060 380
rect 1950 272 1982 318
rect 2028 272 2060 318
rect 1950 210 2060 272
rect 2120 210 2170 380
rect 2230 318 2340 380
rect 2230 272 2262 318
rect 2308 272 2340 318
rect 2230 210 2340 272
rect 2400 318 2500 380
rect 2400 272 2432 318
rect 2478 272 2500 318
rect 2400 210 2500 272
rect 2590 318 2690 380
rect 2590 272 2612 318
rect 2658 272 2690 318
rect 2590 210 2690 272
rect 2750 210 2800 380
rect 2860 318 2970 380
rect 2860 272 2892 318
rect 2938 272 2970 318
rect 2860 210 2970 272
rect 3030 318 3130 380
rect 3030 272 3062 318
rect 3108 272 3130 318
rect 3030 210 3130 272
rect 3220 318 3320 380
rect 3220 272 3242 318
rect 3288 272 3320 318
rect 3220 210 3320 272
rect 3380 318 3490 380
rect 3380 272 3412 318
rect 3458 272 3490 318
rect 3380 210 3490 272
rect 3550 318 3650 380
rect 3550 272 3582 318
rect 3628 272 3650 318
rect 3550 210 3650 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 350 1450
rect 250 1163 282 1397
rect 328 1163 350 1397
rect 250 1110 350 1163
rect 410 1397 510 1450
rect 410 1163 432 1397
rect 478 1163 510 1397
rect 410 1110 510 1163
rect 570 1425 680 1450
rect 570 1285 602 1425
rect 648 1285 680 1425
rect 570 1110 680 1285
rect 740 1425 850 1450
rect 740 1285 772 1425
rect 818 1285 850 1425
rect 740 1110 850 1285
rect 910 1425 1010 1450
rect 910 1285 942 1425
rect 988 1285 1010 1425
rect 910 1110 1010 1285
rect 1070 1397 1170 1450
rect 1070 1163 1092 1397
rect 1138 1163 1170 1397
rect 1070 1110 1170 1163
rect 1230 1110 1330 1450
rect 1390 1397 1500 1450
rect 1390 1163 1422 1397
rect 1468 1163 1500 1397
rect 1390 1110 1500 1163
rect 1560 1110 1610 1450
rect 1670 1397 1780 1450
rect 1670 1163 1702 1397
rect 1748 1163 1780 1397
rect 1670 1110 1780 1163
rect 1840 1110 1890 1450
rect 1950 1425 2060 1450
rect 1950 1285 1982 1425
rect 2028 1285 2060 1425
rect 1950 1110 2060 1285
rect 2120 1110 2170 1450
rect 2230 1425 2340 1450
rect 2230 1285 2262 1425
rect 2308 1285 2340 1425
rect 2230 1110 2340 1285
rect 2400 1397 2500 1450
rect 2400 1163 2432 1397
rect 2478 1163 2500 1397
rect 2400 1110 2500 1163
rect 2560 1430 2660 1450
rect 2560 1290 2582 1430
rect 2628 1290 2660 1430
rect 2560 1110 2660 1290
rect 2720 1428 2830 1450
rect 2720 1382 2752 1428
rect 2798 1382 2830 1428
rect 2720 1110 2830 1382
rect 2890 1388 3000 1450
rect 2890 1342 2922 1388
rect 2968 1342 3000 1388
rect 2890 1110 3000 1342
rect 3060 1397 3160 1450
rect 3060 1163 3092 1397
rect 3138 1163 3160 1397
rect 3060 1110 3160 1163
rect 3220 1397 3320 1450
rect 3220 1163 3242 1397
rect 3288 1163 3320 1397
rect 3220 1110 3320 1163
rect 3380 1397 3490 1450
rect 3380 1163 3412 1397
rect 3458 1163 3490 1397
rect 3380 1110 3490 1163
rect 3550 1397 3650 1450
rect 3550 1163 3582 1397
rect 3628 1163 3650 1397
rect 3550 1110 3650 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 462 272 508 318
rect 632 272 678 318
rect 912 272 958 318
rect 1092 272 1138 318
rect 1422 272 1468 318
rect 1702 232 1748 278
rect 1982 272 2028 318
rect 2262 272 2308 318
rect 2432 272 2478 318
rect 2612 272 2658 318
rect 2892 272 2938 318
rect 3062 272 3108 318
rect 3242 272 3288 318
rect 3412 272 3458 318
rect 3582 272 3628 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 432 1163 478 1397
rect 602 1285 648 1425
rect 772 1285 818 1425
rect 942 1285 988 1425
rect 1092 1163 1138 1397
rect 1422 1163 1468 1397
rect 1702 1163 1748 1397
rect 1982 1285 2028 1425
rect 2262 1285 2308 1425
rect 2432 1163 2478 1397
rect 2582 1290 2628 1430
rect 2752 1382 2798 1428
rect 2922 1342 2968 1388
rect 3092 1163 3138 1397
rect 3242 1163 3288 1397
rect 3412 1163 3458 1397
rect 3582 1163 3628 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 550 118 700 140
rect 550 72 602 118
rect 648 72 700 118
rect 550 50 700 72
rect 790 118 940 140
rect 790 72 842 118
rect 888 72 940 118
rect 790 50 940 72
rect 1030 118 1180 140
rect 1030 72 1082 118
rect 1128 72 1180 118
rect 1030 50 1180 72
rect 1270 118 1420 140
rect 1270 72 1322 118
rect 1368 72 1420 118
rect 1270 50 1420 72
rect 1510 118 1660 140
rect 1510 72 1562 118
rect 1608 72 1660 118
rect 1510 50 1660 72
rect 1750 118 1900 140
rect 1750 72 1802 118
rect 1848 72 1900 118
rect 1750 50 1900 72
rect 1990 118 2140 140
rect 1990 72 2042 118
rect 2088 72 2140 118
rect 1990 50 2140 72
rect 2230 118 2380 140
rect 2230 72 2282 118
rect 2328 72 2380 118
rect 2230 50 2380 72
rect 2470 118 2620 140
rect 2470 72 2522 118
rect 2568 72 2620 118
rect 2470 50 2620 72
rect 2710 118 2860 140
rect 2710 72 2762 118
rect 2808 72 2860 118
rect 2710 50 2860 72
rect 2950 118 3100 140
rect 2950 72 3002 118
rect 3048 72 3100 118
rect 2950 50 3100 72
rect 3190 118 3340 140
rect 3190 72 3242 118
rect 3288 72 3340 118
rect 3190 50 3340 72
rect 3430 118 3580 140
rect 3430 72 3482 118
rect 3528 72 3580 118
rect 3430 50 3580 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 310 1588 460 1610
rect 310 1542 362 1588
rect 408 1542 460 1588
rect 310 1520 460 1542
rect 550 1588 700 1610
rect 550 1542 602 1588
rect 648 1542 700 1588
rect 550 1520 700 1542
rect 790 1588 940 1610
rect 790 1542 842 1588
rect 888 1542 940 1588
rect 790 1520 940 1542
rect 1030 1588 1180 1610
rect 1030 1542 1082 1588
rect 1128 1542 1180 1588
rect 1030 1520 1180 1542
rect 1270 1588 1420 1610
rect 1270 1542 1322 1588
rect 1368 1542 1420 1588
rect 1270 1520 1420 1542
rect 1510 1588 1660 1610
rect 1510 1542 1562 1588
rect 1608 1542 1660 1588
rect 1510 1520 1660 1542
rect 1750 1588 1900 1610
rect 1750 1542 1802 1588
rect 1848 1542 1900 1588
rect 1750 1520 1900 1542
rect 1990 1588 2140 1610
rect 1990 1542 2042 1588
rect 2088 1542 2140 1588
rect 1990 1520 2140 1542
rect 2230 1588 2380 1610
rect 2230 1542 2282 1588
rect 2328 1542 2380 1588
rect 2230 1520 2380 1542
rect 2470 1588 2620 1610
rect 2470 1542 2522 1588
rect 2568 1542 2620 1588
rect 2470 1520 2620 1542
rect 2710 1588 2860 1610
rect 2710 1542 2762 1588
rect 2808 1542 2860 1588
rect 2710 1520 2860 1542
rect 2950 1588 3100 1610
rect 2950 1542 3002 1588
rect 3048 1542 3100 1588
rect 2950 1520 3100 1542
rect 3190 1588 3340 1610
rect 3190 1542 3242 1588
rect 3288 1542 3340 1588
rect 3190 1520 3340 1542
rect 3430 1588 3580 1610
rect 3430 1542 3482 1588
rect 3528 1542 3580 1588
rect 3430 1520 3580 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 602 72 648 118
rect 842 72 888 118
rect 1082 72 1128 118
rect 1322 72 1368 118
rect 1562 72 1608 118
rect 1802 72 1848 118
rect 2042 72 2088 118
rect 2282 72 2328 118
rect 2522 72 2568 118
rect 2762 72 2808 118
rect 3002 72 3048 118
rect 3242 72 3288 118
rect 3482 72 3528 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 362 1542 408 1588
rect 602 1542 648 1588
rect 842 1542 888 1588
rect 1082 1542 1128 1588
rect 1322 1542 1368 1588
rect 1562 1542 1608 1588
rect 1802 1542 1848 1588
rect 2042 1542 2088 1588
rect 2282 1542 2328 1588
rect 2522 1542 2568 1588
rect 2762 1542 2808 1588
rect 3002 1542 3048 1588
rect 3242 1542 3288 1588
rect 3482 1542 3528 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 510 1450 570 1500
rect 680 1450 740 1500
rect 850 1450 910 1500
rect 1170 1450 1230 1500
rect 1330 1450 1390 1500
rect 1500 1450 1560 1500
rect 1610 1450 1670 1500
rect 1780 1450 1840 1500
rect 1890 1450 1950 1500
rect 2060 1450 2120 1500
rect 2170 1450 2230 1500
rect 2340 1450 2400 1500
rect 2660 1450 2720 1500
rect 2830 1450 2890 1500
rect 3000 1450 3060 1500
rect 3320 1450 3380 1500
rect 3490 1450 3550 1500
rect 190 1060 250 1110
rect 120 1038 250 1060
rect 120 992 142 1038
rect 188 992 250 1038
rect 120 970 250 992
rect 190 380 250 970
rect 510 800 570 1110
rect 680 930 740 1110
rect 680 903 800 930
rect 680 857 707 903
rect 753 857 800 903
rect 680 830 800 857
rect 510 773 630 800
rect 510 727 557 773
rect 603 727 630 773
rect 510 700 630 727
rect 510 650 570 700
rect 510 610 600 650
rect 540 380 600 610
rect 680 470 740 830
rect 850 800 910 1110
rect 1170 800 1230 1110
rect 1330 930 1390 1110
rect 1330 903 1430 930
rect 1330 857 1357 903
rect 1403 857 1430 903
rect 1330 830 1430 857
rect 850 773 990 800
rect 850 727 907 773
rect 953 727 990 773
rect 850 700 990 727
rect 1170 773 1290 800
rect 1170 727 1217 773
rect 1263 727 1290 773
rect 1170 700 1290 727
rect 850 470 910 700
rect 680 430 770 470
rect 710 380 770 430
rect 820 430 910 470
rect 820 380 880 430
rect 1170 380 1230 700
rect 1500 660 1560 1110
rect 1610 1060 1670 1110
rect 1780 1060 1840 1110
rect 1610 1033 1840 1060
rect 1610 990 1647 1033
rect 1620 987 1647 990
rect 1693 990 1840 1033
rect 1693 987 1720 990
rect 1620 940 1720 987
rect 1890 660 1950 1110
rect 2060 930 2120 1110
rect 2020 903 2120 930
rect 2020 857 2047 903
rect 2093 857 2120 903
rect 2020 830 2120 857
rect 2170 800 2230 1110
rect 2340 930 2400 1110
rect 2340 903 2440 930
rect 2340 857 2367 903
rect 2413 857 2440 903
rect 2340 830 2440 857
rect 2160 773 2260 800
rect 2160 727 2187 773
rect 2233 727 2260 773
rect 2160 700 2260 727
rect 2020 660 2120 670
rect 1330 643 2120 660
rect 1330 600 2047 643
rect 1330 380 1390 600
rect 2020 597 2047 600
rect 2093 597 2120 643
rect 2020 570 2120 597
rect 1460 513 1560 540
rect 1620 520 1720 540
rect 1460 467 1487 513
rect 1533 467 1560 513
rect 1460 440 1560 467
rect 1500 380 1560 440
rect 1610 513 1840 520
rect 1610 467 1647 513
rect 1693 467 1840 513
rect 1610 440 1840 467
rect 1610 380 1670 440
rect 1780 380 1840 440
rect 1890 503 1990 530
rect 1890 457 1917 503
rect 1963 457 1990 503
rect 1890 430 1990 457
rect 1890 380 1950 430
rect 2060 380 2120 570
rect 2170 380 2230 700
rect 2340 380 2400 830
rect 2660 530 2720 1110
rect 2830 930 2890 1110
rect 2770 903 2890 930
rect 2770 857 2817 903
rect 2863 857 2890 903
rect 2770 830 2890 857
rect 2580 503 2720 530
rect 2580 457 2617 503
rect 2663 470 2720 503
rect 2830 470 2890 830
rect 3000 650 3060 1110
rect 3320 670 3380 1110
rect 3490 930 3550 1110
rect 3430 903 3550 930
rect 3430 857 3457 903
rect 3503 857 3550 903
rect 3430 830 3550 857
rect 2663 457 2750 470
rect 2580 430 2750 457
rect 2690 380 2750 430
rect 2800 430 2890 470
rect 2970 610 3060 650
rect 3260 643 3380 670
rect 2970 530 3030 610
rect 3260 597 3307 643
rect 3353 597 3380 643
rect 3260 570 3380 597
rect 2970 503 3090 530
rect 2970 457 3017 503
rect 3063 457 3090 503
rect 2970 430 3090 457
rect 2800 380 2860 430
rect 2970 380 3030 430
rect 3320 380 3380 570
rect 3490 380 3550 830
rect 190 160 250 210
rect 540 160 600 210
rect 710 160 770 210
rect 820 160 880 210
rect 1170 160 1230 210
rect 1330 160 1390 210
rect 1500 160 1560 210
rect 1610 160 1670 210
rect 1780 160 1840 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2170 160 2230 210
rect 2340 160 2400 210
rect 2690 160 2750 210
rect 2800 160 2860 210
rect 2970 160 3030 210
rect 3320 160 3380 210
rect 3490 160 3550 210
<< polycontact >>
rect 142 992 188 1038
rect 707 857 753 903
rect 557 727 603 773
rect 1357 857 1403 903
rect 907 727 953 773
rect 1217 727 1263 773
rect 1647 987 1693 1033
rect 2047 857 2093 903
rect 2367 857 2413 903
rect 2187 727 2233 773
rect 2047 597 2093 643
rect 1487 467 1533 513
rect 1647 467 1693 513
rect 1917 457 1963 503
rect 2817 857 2863 903
rect 2617 457 2663 503
rect 3457 857 3503 903
rect 3307 597 3353 643
rect 3017 457 3063 503
<< metal1 >>
rect 0 1588 3740 1660
rect 0 1542 112 1588
rect 158 1542 362 1588
rect 408 1542 602 1588
rect 648 1542 842 1588
rect 888 1542 1082 1588
rect 1128 1542 1322 1588
rect 1368 1542 1562 1588
rect 1608 1542 1802 1588
rect 1848 1542 2042 1588
rect 2088 1542 2282 1588
rect 2328 1542 2522 1588
rect 2568 1542 2762 1588
rect 2808 1542 3002 1588
rect 3048 1542 3242 1588
rect 3288 1542 3482 1588
rect 3528 1542 3740 1588
rect 0 1520 3740 1542
rect 110 1397 160 1520
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1110 160 1163
rect 280 1397 330 1450
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 110 1038 210 1040
rect 110 1036 142 1038
rect 110 984 134 1036
rect 188 992 210 1038
rect 186 984 210 992
rect 110 980 210 984
rect 280 520 330 1163
rect 430 1397 480 1450
rect 430 1163 432 1397
rect 478 1163 480 1397
rect 430 570 480 1163
rect 600 1425 650 1450
rect 600 1285 602 1425
rect 648 1285 650 1425
rect 600 1210 650 1285
rect 770 1425 820 1520
rect 770 1285 772 1425
rect 818 1285 820 1425
rect 770 1260 820 1285
rect 940 1425 990 1450
rect 940 1285 942 1425
rect 988 1285 990 1425
rect 940 1210 990 1285
rect 600 1160 990 1210
rect 1090 1397 1140 1520
rect 1090 1163 1092 1397
rect 1138 1163 1140 1397
rect 1090 1110 1140 1163
rect 1420 1397 1470 1450
rect 1420 1163 1422 1397
rect 1468 1163 1470 1397
rect 1420 1060 1470 1163
rect 1700 1397 1750 1520
rect 1700 1163 1702 1397
rect 1748 1163 1750 1397
rect 1980 1425 2030 1450
rect 1980 1285 1982 1425
rect 2028 1285 2030 1425
rect 1980 1260 2030 1285
rect 2260 1425 2310 1520
rect 2260 1285 2262 1425
rect 2308 1285 2310 1425
rect 2260 1260 2310 1285
rect 2430 1397 2480 1450
rect 1700 1110 1750 1163
rect 1800 1210 2030 1260
rect 1090 1010 1470 1060
rect 1620 1033 1720 1040
rect 680 906 780 910
rect 680 854 704 906
rect 756 854 780 906
rect 680 850 780 854
rect 1090 780 1140 1010
rect 1620 987 1647 1033
rect 1693 987 1720 1033
rect 1620 980 1720 987
rect 1330 906 1560 910
rect 1330 903 1484 906
rect 1330 857 1357 903
rect 1403 857 1484 903
rect 1330 854 1484 857
rect 1536 854 1560 906
rect 1330 850 1560 854
rect 530 776 630 780
rect 530 724 554 776
rect 606 724 630 776
rect 530 720 630 724
rect 880 776 1140 780
rect 880 724 904 776
rect 956 724 1140 776
rect 880 720 1140 724
rect 1190 776 1290 780
rect 1190 724 1214 776
rect 1266 724 1290 776
rect 1190 720 1290 724
rect 430 520 680 570
rect 900 520 950 530
rect 1090 520 1140 720
rect 1480 520 1540 850
rect 1640 520 1700 980
rect 1800 760 1850 1210
rect 2430 1163 2432 1397
rect 2478 1163 2480 1397
rect 2580 1430 2630 1450
rect 2580 1290 2582 1430
rect 2628 1310 2630 1430
rect 2750 1428 2800 1520
rect 2750 1382 2752 1428
rect 2798 1382 2800 1428
rect 2750 1360 2800 1382
rect 2920 1388 2970 1450
rect 2920 1342 2922 1388
rect 2968 1342 2970 1388
rect 2920 1310 2970 1342
rect 2628 1290 2970 1310
rect 2580 1260 2970 1290
rect 3090 1397 3140 1450
rect 2150 1036 2250 1040
rect 2150 984 2174 1036
rect 2226 984 2250 1036
rect 2150 980 2250 984
rect 2430 1020 2480 1163
rect 3090 1163 3092 1397
rect 3138 1163 3140 1397
rect 2610 1040 2670 1060
rect 3090 1040 3140 1163
rect 3240 1397 3290 1450
rect 3240 1163 3242 1397
rect 3288 1163 3290 1397
rect 2610 1036 3170 1040
rect 1790 710 1850 760
rect 1910 906 2120 910
rect 1910 854 2044 906
rect 2096 854 2120 906
rect 1910 850 2120 854
rect 260 516 360 520
rect 260 464 284 516
rect 336 464 360 516
rect 260 460 360 464
rect 630 516 980 520
rect 630 464 904 516
rect 956 464 980 516
rect 1090 470 1290 520
rect 630 460 980 464
rect 280 450 340 460
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 450
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 460 318 510 380
rect 460 272 462 318
rect 508 272 510 318
rect 460 140 510 272
rect 630 318 680 460
rect 900 450 950 460
rect 1210 380 1290 470
rect 1460 513 1560 520
rect 1460 467 1487 513
rect 1533 467 1560 513
rect 1460 460 1560 467
rect 1620 516 1720 520
rect 1620 464 1644 516
rect 1696 464 1720 516
rect 1620 460 1720 464
rect 1790 390 1840 710
rect 1910 510 1970 850
rect 2170 780 2230 980
rect 2430 970 2540 1020
rect 2340 906 2440 910
rect 2340 854 2364 906
rect 2416 854 2440 906
rect 2340 850 2440 854
rect 2490 780 2540 970
rect 2610 984 2614 1036
rect 2666 984 3094 1036
rect 3146 984 3170 1036
rect 2610 980 3170 984
rect 2610 960 2670 980
rect 2790 906 2890 910
rect 2790 854 2814 906
rect 2866 854 2890 906
rect 2790 850 2890 854
rect 2160 776 2260 780
rect 2160 724 2184 776
rect 2236 724 2260 776
rect 2160 720 2260 724
rect 2430 730 2540 780
rect 2020 646 2120 650
rect 2020 594 2044 646
rect 2096 594 2120 646
rect 2020 590 2120 594
rect 2430 646 2490 730
rect 3090 650 3140 980
rect 3240 910 3290 1163
rect 3410 1397 3460 1520
rect 3410 1163 3412 1397
rect 3458 1163 3460 1397
rect 3410 1110 3460 1163
rect 3580 1397 3630 1450
rect 3580 1163 3582 1397
rect 3628 1163 3630 1397
rect 3580 1050 3630 1163
rect 3580 1036 3680 1050
rect 3580 984 3604 1036
rect 3656 984 3680 1036
rect 3580 980 3680 984
rect 3580 970 3670 980
rect 3240 906 3530 910
rect 3240 854 3454 906
rect 3506 854 3530 906
rect 3240 850 3530 854
rect 2430 594 2434 646
rect 2486 594 2490 646
rect 2430 570 2490 594
rect 2890 646 3380 650
rect 2890 594 3304 646
rect 3356 594 3380 646
rect 2890 590 3380 594
rect 1890 503 1990 510
rect 1890 457 1917 503
rect 1963 457 1990 503
rect 1890 450 1990 457
rect 1790 386 2060 390
rect 630 272 632 318
rect 678 272 680 318
rect 630 210 680 272
rect 910 318 960 380
rect 910 272 912 318
rect 958 272 960 318
rect 910 140 960 272
rect 1090 318 1140 380
rect 1210 330 1470 380
rect 1790 340 1984 386
rect 1090 272 1092 318
rect 1138 272 1140 318
rect 1090 140 1140 272
rect 1420 318 1470 330
rect 1420 272 1422 318
rect 1468 272 1470 318
rect 1980 334 1984 340
rect 2036 334 2060 386
rect 1980 330 2060 334
rect 1980 318 2030 330
rect 1420 210 1470 272
rect 1700 278 1750 300
rect 1700 232 1702 278
rect 1748 232 1750 278
rect 1700 140 1750 232
rect 1980 272 1982 318
rect 2028 272 2030 318
rect 1980 210 2030 272
rect 2260 318 2310 380
rect 2260 272 2262 318
rect 2308 272 2310 318
rect 2260 140 2310 272
rect 2430 318 2480 570
rect 2590 506 2690 510
rect 2590 454 2614 506
rect 2666 454 2690 506
rect 2590 450 2690 454
rect 2430 272 2432 318
rect 2478 272 2480 318
rect 2430 210 2480 272
rect 2610 318 2660 380
rect 2610 272 2612 318
rect 2658 272 2660 318
rect 2610 140 2660 272
rect 2890 318 2940 590
rect 2990 506 3090 510
rect 2990 454 3014 506
rect 3066 454 3090 506
rect 3460 480 3510 850
rect 2990 450 3090 454
rect 3240 430 3510 480
rect 2890 272 2892 318
rect 2938 272 2940 318
rect 2890 210 2940 272
rect 3060 318 3110 380
rect 3060 272 3062 318
rect 3108 272 3110 318
rect 3060 140 3110 272
rect 3240 318 3290 430
rect 3240 272 3242 318
rect 3288 272 3290 318
rect 3240 210 3290 272
rect 3410 318 3460 380
rect 3410 272 3412 318
rect 3458 272 3460 318
rect 3410 140 3460 272
rect 3580 318 3630 970
rect 3580 272 3582 318
rect 3628 272 3630 318
rect 3580 210 3630 272
rect 0 118 3740 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 602 118
rect 648 72 842 118
rect 888 72 1082 118
rect 1128 72 1322 118
rect 1368 72 1562 118
rect 1608 72 1802 118
rect 1848 72 2042 118
rect 2088 72 2282 118
rect 2328 72 2522 118
rect 2568 72 2762 118
rect 2808 72 3002 118
rect 3048 72 3242 118
rect 3288 72 3482 118
rect 3528 72 3740 118
rect 0 0 3740 72
<< via1 >>
rect 134 992 142 1036
rect 142 992 186 1036
rect 134 984 186 992
rect 704 903 756 906
rect 704 857 707 903
rect 707 857 753 903
rect 753 857 756 903
rect 704 854 756 857
rect 1484 854 1536 906
rect 554 773 606 776
rect 554 727 557 773
rect 557 727 603 773
rect 603 727 606 773
rect 554 724 606 727
rect 904 773 956 776
rect 904 727 907 773
rect 907 727 953 773
rect 953 727 956 773
rect 904 724 956 727
rect 1214 773 1266 776
rect 1214 727 1217 773
rect 1217 727 1263 773
rect 1263 727 1266 773
rect 1214 724 1266 727
rect 2174 984 2226 1036
rect 2044 903 2096 906
rect 2044 857 2047 903
rect 2047 857 2093 903
rect 2093 857 2096 903
rect 2044 854 2096 857
rect 284 464 336 516
rect 904 464 956 516
rect 1644 513 1696 516
rect 1644 467 1647 513
rect 1647 467 1693 513
rect 1693 467 1696 513
rect 1644 464 1696 467
rect 2364 903 2416 906
rect 2364 857 2367 903
rect 2367 857 2413 903
rect 2413 857 2416 903
rect 2364 854 2416 857
rect 2614 984 2666 1036
rect 3094 984 3146 1036
rect 2814 903 2866 906
rect 2814 857 2817 903
rect 2817 857 2863 903
rect 2863 857 2866 903
rect 2814 854 2866 857
rect 2184 773 2236 776
rect 2184 727 2187 773
rect 2187 727 2233 773
rect 2233 727 2236 773
rect 2184 724 2236 727
rect 2044 643 2096 646
rect 2044 597 2047 643
rect 2047 597 2093 643
rect 2093 597 2096 643
rect 2044 594 2096 597
rect 3604 984 3656 1036
rect 3454 903 3506 906
rect 3454 857 3457 903
rect 3457 857 3503 903
rect 3503 857 3506 903
rect 3454 854 3506 857
rect 2434 594 2486 646
rect 3304 643 3356 646
rect 3304 597 3307 643
rect 3307 597 3353 643
rect 3353 597 3356 643
rect 3304 594 3356 597
rect 1984 334 2036 386
rect 2614 503 2666 506
rect 2614 457 2617 503
rect 2617 457 2663 503
rect 2663 457 2666 503
rect 2614 454 2666 457
rect 3014 503 3066 506
rect 3014 457 3017 503
rect 3017 457 3063 503
rect 3063 457 3066 503
rect 3014 454 3066 457
<< metal2 >>
rect 700 1110 2870 1170
rect 110 1036 210 1050
rect 110 984 134 1036
rect 186 984 210 1036
rect 110 970 210 984
rect 700 920 760 1110
rect 2160 1040 2240 1050
rect 2600 1040 2680 1050
rect 2150 1036 2690 1040
rect 2150 984 2174 1036
rect 2226 984 2614 1036
rect 2666 984 2690 1036
rect 2150 980 2690 984
rect 2160 970 2240 980
rect 2600 970 2680 980
rect 2810 920 2870 1110
rect 3070 1036 3170 1050
rect 3590 1040 3670 1050
rect 3070 984 3094 1036
rect 3146 984 3170 1036
rect 3070 970 3170 984
rect 3580 1036 3680 1040
rect 3580 984 3604 1036
rect 3656 984 3680 1036
rect 3580 980 3680 984
rect 3590 970 3670 980
rect 680 906 780 920
rect 680 854 704 906
rect 756 854 780 906
rect 680 840 780 854
rect 1460 910 1550 920
rect 2020 910 2120 920
rect 2350 910 2430 920
rect 1460 906 2440 910
rect 1460 854 1484 906
rect 1536 854 2044 906
rect 2096 854 2364 906
rect 2416 854 2440 906
rect 1460 850 2440 854
rect 2790 906 2890 920
rect 3440 910 3520 920
rect 2790 854 2814 906
rect 2866 854 2890 906
rect 1460 840 1550 850
rect 2020 840 2120 850
rect 2350 840 2430 850
rect 2790 840 2890 854
rect 3430 906 3530 910
rect 3430 854 3454 906
rect 3506 854 3530 906
rect 3430 850 3530 854
rect 3440 840 3520 850
rect 530 776 630 790
rect 530 724 554 776
rect 606 724 630 776
rect 530 710 630 724
rect 880 776 980 790
rect 880 724 904 776
rect 956 724 980 776
rect 880 710 980 724
rect 1190 776 1290 790
rect 2170 780 2250 790
rect 1190 724 1214 776
rect 1266 724 1290 776
rect 1190 710 1290 724
rect 2160 776 2260 780
rect 2160 724 2184 776
rect 2236 724 2260 776
rect 2160 720 2260 724
rect 2170 710 2250 720
rect 260 520 360 530
rect 550 520 610 710
rect 2030 650 2110 660
rect 2420 650 2500 660
rect 3290 650 3370 660
rect 2020 646 2520 650
rect 2020 594 2044 646
rect 2096 594 2434 646
rect 2486 594 2520 646
rect 2020 590 2520 594
rect 3220 646 3380 650
rect 3220 594 3304 646
rect 3356 594 3380 646
rect 3220 590 3380 594
rect 2030 580 2110 590
rect 2420 580 2500 590
rect 3290 580 3370 590
rect 260 516 610 520
rect 260 464 284 516
rect 336 464 610 516
rect 260 460 610 464
rect 260 450 360 460
rect 550 260 610 460
rect 880 520 980 530
rect 1630 520 1710 530
rect 880 516 1720 520
rect 880 464 904 516
rect 956 464 1644 516
rect 1696 464 1720 516
rect 880 460 1720 464
rect 2590 506 2690 520
rect 880 450 980 460
rect 1630 450 1710 460
rect 2590 454 2614 506
rect 2666 454 2690 506
rect 2590 440 2690 454
rect 2970 506 3090 520
rect 2970 454 3014 506
rect 3066 454 3090 506
rect 2970 440 3090 454
rect 1970 390 2050 400
rect 2590 390 2670 440
rect 1960 386 2670 390
rect 1960 334 1984 386
rect 2036 334 2670 386
rect 1960 330 2670 334
rect 1970 320 2050 330
rect 2970 260 3030 440
rect 550 200 3030 260
<< labels >>
rlabel via1 s 1214 724 1266 776 4 D
port 1 nsew signal input
rlabel via1 s 3604 984 3656 1036 4 Q
port 2 nsew signal output
rlabel via1 s 3454 854 3506 906 4 QN
port 3 nsew signal output
rlabel via1 s 134 984 186 1036 4 RN
port 4 nsew signal input
rlabel via1 s 2814 854 2866 906 4 SN
port 5 nsew signal output
rlabel via1 s 2364 854 2416 906 4 CLK
port 6 nsew clock input
rlabel metal1 s 110 1110 160 1660 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 770 1260 820 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1090 1110 1140 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1700 1110 1750 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2260 1260 2310 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2750 1360 2800 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3410 1110 3460 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3740 1660 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 460 0 510 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 910 0 960 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1090 0 1140 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1700 0 1750 300 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2260 0 2310 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2610 0 2660 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3060 0 3110 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3410 0 3460 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3740 140 1 VSS
port 8 nsew ground bidirectional abutment
rlabel via1 s 2044 854 2096 906 1 CLK
port 6 nsew clock input
rlabel via1 s 1484 854 1536 906 1 CLK
port 6 nsew clock input
rlabel metal2 s 1460 840 1550 920 1 CLK
port 6 nsew clock input
rlabel metal2 s 2020 840 2120 920 1 CLK
port 6 nsew clock input
rlabel metal2 s 2350 840 2430 920 1 CLK
port 6 nsew clock input
rlabel metal2 s 1460 850 2440 910 1 CLK
port 6 nsew clock input
rlabel metal1 s 1480 460 1540 910 1 CLK
port 6 nsew clock input
rlabel metal1 s 1460 460 1560 520 1 CLK
port 6 nsew clock input
rlabel metal1 s 1330 850 1560 910 1 CLK
port 6 nsew clock input
rlabel metal1 s 1910 450 1970 910 1 CLK
port 6 nsew clock input
rlabel metal1 s 1890 450 1990 510 1 CLK
port 6 nsew clock input
rlabel metal1 s 1910 850 2120 910 1 CLK
port 6 nsew clock input
rlabel metal1 s 2340 850 2440 910 1 CLK
port 6 nsew clock input
rlabel metal2 s 1190 710 1290 790 1 D
port 1 nsew signal input
rlabel metal1 s 1190 720 1290 780 1 D
port 1 nsew signal input
rlabel metal2 s 3590 970 3670 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3580 980 3680 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 3580 210 3630 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 3580 970 3670 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 3580 980 3680 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3440 840 3520 920 1 QN
port 3 nsew signal output
rlabel metal2 s 3430 850 3530 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3240 210 3290 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3240 850 3290 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 3240 430 3510 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3460 430 3510 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3240 850 3530 910 1 QN
port 3 nsew signal output
rlabel metal2 s 110 970 210 1050 1 RN
port 4 nsew signal input
rlabel metal1 s 110 980 210 1040 1 RN
port 4 nsew signal input
rlabel via1 s 704 854 756 906 1 SN
port 5 nsew signal output
rlabel metal2 s 700 840 760 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 680 840 780 920 1 SN
port 5 nsew signal output
rlabel metal2 s 2810 840 2870 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 700 1110 2870 1170 1 SN
port 5 nsew signal output
rlabel metal2 s 2790 840 2890 920 1 SN
port 5 nsew signal output
rlabel metal1 s 680 850 780 910 1 SN
port 5 nsew signal output
rlabel metal1 s 2790 850 2890 910 1 SN
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3740 1660
string GDS_END 344892
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 315458
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
