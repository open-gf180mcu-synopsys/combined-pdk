magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 377 4902 870
rect -86 352 1827 377
rect 3033 352 4902 377
<< pwell >>
rect 1827 352 3033 377
rect -86 -86 4902 352
<< mvnmos >>
rect 124 151 244 232
rect 348 151 468 232
rect 716 156 836 228
rect 940 156 1060 228
rect 1164 156 1284 228
rect 1353 156 1473 228
rect 1577 156 1697 228
rect 1793 156 1913 228
rect 2105 156 2225 228
rect 2329 156 2449 228
rect 2961 151 3081 232
rect 3129 151 3249 232
rect 3397 69 3517 232
rect 3621 69 3741 232
rect 3861 69 3981 232
rect 4085 69 4205 232
rect 4309 69 4429 232
rect 4533 69 4653 232
<< mvpmos >>
rect 144 472 244 645
rect 348 472 448 645
rect 736 527 836 628
rect 940 527 1040 628
rect 1193 527 1293 628
rect 1373 527 1473 628
rect 1689 527 1789 644
rect 1893 527 1993 644
rect 2393 497 2493 580
rect 2597 497 2697 580
rect 2945 504 3045 660
rect 3149 504 3249 660
rect 3417 504 3517 715
rect 3621 504 3721 715
rect 3861 472 3961 715
rect 4105 472 4205 715
rect 4309 472 4409 715
rect 4553 472 4653 715
<< mvndiff >>
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 151 124 173
rect 244 210 348 232
rect 244 164 273 210
rect 319 164 348 210
rect 244 151 348 164
rect 468 219 556 232
rect 1973 244 2045 257
rect 1973 228 1986 244
rect 468 173 497 219
rect 543 173 556 219
rect 468 151 556 173
rect 628 215 716 228
rect 628 169 641 215
rect 687 169 716 215
rect 628 156 716 169
rect 836 215 940 228
rect 836 169 865 215
rect 911 169 940 215
rect 836 156 940 169
rect 1060 215 1164 228
rect 1060 169 1089 215
rect 1135 169 1164 215
rect 1060 156 1164 169
rect 1284 156 1353 228
rect 1473 215 1577 228
rect 1473 169 1502 215
rect 1548 169 1577 215
rect 1473 156 1577 169
rect 1697 156 1793 228
rect 1913 198 1986 228
rect 2032 228 2045 244
rect 2509 244 2581 257
rect 2509 228 2522 244
rect 2032 198 2105 228
rect 1913 156 2105 198
rect 2225 215 2329 228
rect 2225 169 2254 215
rect 2300 169 2329 215
rect 2225 156 2329 169
rect 2449 198 2522 228
rect 2568 198 2581 244
rect 2449 156 2581 198
rect 2829 244 2901 257
rect 2829 198 2842 244
rect 2888 232 2901 244
rect 2888 198 2961 232
rect 2829 151 2961 198
rect 3081 151 3129 232
rect 3249 167 3397 232
rect 3249 151 3322 167
rect 3309 121 3322 151
rect 3368 121 3397 167
rect 3309 69 3397 121
rect 3517 167 3621 232
rect 3517 121 3546 167
rect 3592 121 3621 167
rect 3517 69 3621 121
rect 3741 167 3861 232
rect 3741 121 3770 167
rect 3816 121 3861 167
rect 3741 69 3861 121
rect 3981 167 4085 232
rect 3981 121 4010 167
rect 4056 121 4085 167
rect 3981 69 4085 121
rect 4205 167 4309 232
rect 4205 121 4234 167
rect 4280 121 4309 167
rect 4205 69 4309 121
rect 4429 167 4533 232
rect 4429 121 4458 167
rect 4504 121 4533 167
rect 4429 69 4533 121
rect 4653 167 4741 232
rect 4653 121 4682 167
rect 4728 121 4741 167
rect 4653 69 4741 121
<< mvpdiff >>
rect 56 632 144 645
rect 56 492 69 632
rect 115 492 144 632
rect 56 472 144 492
rect 244 632 348 645
rect 244 586 273 632
rect 319 586 348 632
rect 244 472 348 586
rect 448 632 536 645
rect 448 492 477 632
rect 523 492 536 632
rect 1533 735 1605 748
rect 1533 689 1546 735
rect 1592 689 1605 735
rect 1533 644 1605 689
rect 2053 647 2125 660
rect 2053 644 2066 647
rect 1533 628 1689 644
rect 646 615 736 628
rect 646 569 659 615
rect 705 569 736 615
rect 646 527 736 569
rect 836 586 940 628
rect 836 540 865 586
rect 911 540 940 586
rect 836 527 940 540
rect 1040 586 1193 628
rect 1040 540 1069 586
rect 1115 540 1193 586
rect 1040 527 1193 540
rect 1293 527 1373 628
rect 1473 527 1689 628
rect 1789 586 1893 644
rect 1789 540 1818 586
rect 1864 540 1893 586
rect 1789 527 1893 540
rect 1993 601 2066 644
rect 2112 601 2125 647
rect 1993 527 2125 601
rect 3317 665 3417 715
rect 3317 660 3341 665
rect 2857 647 2945 660
rect 2857 601 2870 647
rect 2916 601 2945 647
rect 2259 556 2393 580
rect 448 472 536 492
rect 2259 510 2272 556
rect 2318 510 2393 556
rect 2259 497 2393 510
rect 2493 556 2597 580
rect 2493 510 2522 556
rect 2568 510 2597 556
rect 2493 497 2597 510
rect 2697 556 2785 580
rect 2697 510 2726 556
rect 2772 510 2785 556
rect 2697 497 2785 510
rect 2857 504 2945 601
rect 3045 566 3149 660
rect 3045 520 3074 566
rect 3120 520 3149 566
rect 3045 504 3149 520
rect 3249 520 3341 660
rect 3387 520 3417 665
rect 3249 504 3417 520
rect 3517 665 3621 715
rect 3517 520 3546 665
rect 3592 520 3621 665
rect 3517 504 3621 520
rect 3721 665 3861 715
rect 3721 520 3750 665
rect 3796 520 3861 665
rect 3721 504 3861 520
rect 3781 472 3861 504
rect 3961 665 4105 715
rect 3961 520 4010 665
rect 4056 520 4105 665
rect 3961 472 4105 520
rect 4205 665 4309 715
rect 4205 520 4234 665
rect 4280 520 4309 665
rect 4205 472 4309 520
rect 4409 665 4553 715
rect 4409 520 4458 665
rect 4504 520 4553 665
rect 4409 472 4553 520
rect 4653 665 4741 715
rect 4653 520 4682 665
rect 4728 520 4741 665
rect 4653 472 4741 520
<< mvndiffc >>
rect 49 173 95 219
rect 273 164 319 210
rect 497 173 543 219
rect 641 169 687 215
rect 865 169 911 215
rect 1089 169 1135 215
rect 1502 169 1548 215
rect 1986 198 2032 244
rect 2254 169 2300 215
rect 2522 198 2568 244
rect 2842 198 2888 244
rect 3322 121 3368 167
rect 3546 121 3592 167
rect 3770 121 3816 167
rect 4010 121 4056 167
rect 4234 121 4280 167
rect 4458 121 4504 167
rect 4682 121 4728 167
<< mvpdiffc >>
rect 69 492 115 632
rect 273 586 319 632
rect 477 492 523 632
rect 1546 689 1592 735
rect 659 569 705 615
rect 865 540 911 586
rect 1069 540 1115 586
rect 1818 540 1864 586
rect 2066 601 2112 647
rect 2870 601 2916 647
rect 2272 510 2318 556
rect 2522 510 2568 556
rect 2726 510 2772 556
rect 3074 520 3120 566
rect 3341 520 3387 665
rect 3546 520 3592 665
rect 3750 520 3796 665
rect 4010 520 4056 665
rect 4234 520 4280 665
rect 4458 520 4504 665
rect 4682 520 4728 665
<< polysilicon >>
rect 348 720 1293 760
rect 144 645 244 690
rect 348 645 448 720
rect 736 628 836 672
rect 940 628 1040 672
rect 1193 628 1293 720
rect 1373 628 1473 672
rect 1893 720 3045 760
rect 1689 644 1789 688
rect 1893 644 1993 720
rect 2393 659 2493 672
rect 2945 660 3045 720
rect 3417 715 3517 760
rect 3621 715 3721 760
rect 3861 715 3961 760
rect 4105 715 4205 760
rect 4309 715 4409 760
rect 4553 715 4653 760
rect 3149 660 3249 704
rect 2393 613 2406 659
rect 2452 613 2493 659
rect 2393 580 2493 613
rect 2597 580 2697 624
rect 144 406 244 472
rect 144 360 157 406
rect 203 360 244 406
rect 144 276 244 360
rect 124 232 244 276
rect 348 336 448 472
rect 348 290 372 336
rect 418 290 448 336
rect 348 276 448 290
rect 736 415 836 527
rect 736 369 749 415
rect 795 369 836 415
rect 736 276 836 369
rect 940 443 1040 527
rect 940 397 977 443
rect 1023 410 1040 443
rect 1193 494 1293 527
rect 1193 448 1234 494
rect 1280 448 1293 494
rect 1193 435 1293 448
rect 1373 491 1473 527
rect 1373 445 1414 491
rect 1460 445 1473 491
rect 1023 397 1147 410
rect 940 351 1147 397
rect 940 324 1284 351
rect 1107 311 1284 324
rect 1164 307 1284 311
rect 348 232 468 276
rect 716 228 836 276
rect 940 228 1060 276
rect 1164 261 1211 307
rect 1257 261 1284 307
rect 1373 276 1473 445
rect 1689 419 1789 527
rect 1893 467 1993 527
rect 1164 228 1284 261
rect 1353 228 1473 276
rect 1577 399 1789 419
rect 1577 353 1590 399
rect 1636 379 1789 399
rect 1636 353 1697 379
rect 1577 228 1697 353
rect 1837 331 1993 467
rect 2393 401 2493 497
rect 1793 327 1993 331
rect 2329 361 2493 401
rect 2597 401 2697 497
rect 2945 415 3045 504
rect 1793 228 1913 327
rect 2105 311 2225 324
rect 2105 265 2162 311
rect 2208 265 2225 311
rect 2105 228 2225 265
rect 2329 228 2449 361
rect 2597 327 2741 401
rect 124 107 244 151
rect 348 64 468 151
rect 716 112 836 156
rect 940 64 1060 156
rect 1164 112 1284 156
rect 1353 112 1473 156
rect 1577 112 1697 156
rect 1793 112 1913 156
rect 348 24 1060 64
rect 2105 64 2225 156
rect 2329 112 2449 156
rect 2641 64 2741 327
rect 2945 369 2958 415
rect 3004 369 3045 415
rect 2945 311 3045 369
rect 2961 301 3045 311
rect 3149 419 3249 504
rect 3149 373 3162 419
rect 3208 373 3249 419
rect 2961 232 3081 301
rect 3149 288 3249 373
rect 3417 351 3517 504
rect 3621 351 3721 504
rect 3861 370 3961 472
rect 4105 370 4205 472
rect 4309 370 4409 472
rect 4553 370 4653 472
rect 3861 357 4653 370
rect 3129 232 3249 288
rect 3397 326 3741 351
rect 3397 280 3410 326
rect 3456 311 3741 326
rect 3456 280 3517 311
rect 3397 232 3517 280
rect 3621 232 3741 311
rect 3861 311 3880 357
rect 4302 311 4653 357
rect 3861 298 4653 311
rect 3861 232 3981 298
rect 4085 232 4205 298
rect 4309 232 4429 298
rect 4533 232 4653 298
rect 2961 107 3081 151
rect 3129 107 3249 151
rect 2105 24 2741 64
rect 3397 24 3517 69
rect 3621 24 3741 69
rect 3861 24 3981 69
rect 4085 24 4205 69
rect 4309 24 4429 69
rect 4533 24 4653 69
<< polycontact >>
rect 2406 613 2452 659
rect 157 360 203 406
rect 372 290 418 336
rect 749 369 795 415
rect 977 397 1023 443
rect 1234 448 1280 494
rect 1414 445 1460 491
rect 1211 261 1257 307
rect 1590 353 1636 399
rect 2162 265 2208 311
rect 2958 369 3004 415
rect 3162 373 3208 419
rect 3410 280 3456 326
rect 3880 311 4302 357
<< metal1 >>
rect 0 735 4816 844
rect 0 724 1546 735
rect 69 632 115 645
rect 262 632 330 724
rect 262 586 273 632
rect 319 586 330 632
rect 477 632 523 645
rect 115 492 418 519
rect 69 472 418 492
rect 56 406 318 426
rect 56 360 157 406
rect 203 360 318 406
rect 56 353 318 360
rect 372 336 418 472
rect 49 290 372 302
rect 49 256 418 290
rect 648 615 716 724
rect 1535 689 1546 724
rect 1592 724 4816 735
rect 1592 689 1603 724
rect 648 569 659 615
rect 705 569 716 615
rect 762 632 1023 678
rect 1654 643 1983 678
rect 762 523 808 632
rect 523 492 808 523
rect 477 476 808 492
rect 854 540 865 586
rect 911 540 922 586
rect 49 219 95 256
rect 477 230 524 476
rect 578 415 806 430
rect 578 369 749 415
rect 795 369 806 415
rect 578 354 806 369
rect 477 219 543 230
rect 49 162 95 173
rect 262 164 273 210
rect 319 164 330 210
rect 262 60 330 164
rect 477 173 497 219
rect 854 215 922 540
rect 977 443 1023 632
rect 1223 632 1983 643
rect 1223 597 1700 632
rect 977 386 1023 397
rect 1069 586 1115 597
rect 1069 399 1115 540
rect 1223 494 1291 597
rect 1223 448 1234 494
rect 1280 448 1291 494
rect 1807 540 1818 586
rect 1864 540 1875 586
rect 1807 491 1875 540
rect 1937 555 1983 632
rect 2055 647 2123 724
rect 2055 601 2066 647
rect 2112 601 2123 647
rect 2169 613 2406 659
rect 2452 613 2463 659
rect 2859 647 2927 724
rect 2169 555 2215 613
rect 2859 601 2870 647
rect 2916 601 2927 647
rect 3341 665 3387 724
rect 2726 556 2772 569
rect 1937 508 2215 555
rect 2261 510 2272 556
rect 2318 510 2329 556
rect 1403 445 1414 491
rect 1460 462 1875 491
rect 2261 462 2329 510
rect 1460 445 2329 462
rect 1807 416 2329 445
rect 2386 510 2522 556
rect 2568 510 2579 556
rect 3074 566 3120 577
rect 2772 520 3074 555
rect 2772 510 3120 520
rect 477 162 543 173
rect 630 169 641 215
rect 687 169 698 215
rect 630 60 698 169
rect 854 169 865 215
rect 911 169 922 215
rect 854 158 922 169
rect 1069 353 1590 399
rect 1636 353 1647 399
rect 1069 215 1135 353
rect 1200 261 1211 307
rect 1257 261 1668 307
rect 1069 169 1089 215
rect 1069 158 1135 169
rect 1491 169 1502 215
rect 1548 169 1559 215
rect 1491 60 1559 169
rect 1622 152 1668 261
rect 1975 244 2043 416
rect 1975 198 1986 244
rect 2032 198 2043 244
rect 2162 311 2208 323
rect 2162 152 2208 265
rect 2386 226 2432 510
rect 2726 508 3120 510
rect 2726 244 2772 508
rect 3341 506 3387 520
rect 3546 665 3592 676
rect 2818 415 3057 430
rect 3546 421 3592 520
rect 3750 665 3796 724
rect 3750 506 3796 520
rect 4010 665 4056 676
rect 2818 369 2958 415
rect 3004 369 3057 415
rect 3151 419 3592 421
rect 3151 373 3162 419
rect 3208 373 3592 419
rect 4010 458 4056 520
rect 4234 665 4280 724
rect 4234 506 4280 520
rect 4334 665 4507 676
rect 4334 520 4458 665
rect 4504 520 4507 665
rect 4334 458 4507 520
rect 4682 665 4728 724
rect 4682 506 4728 520
rect 4010 412 4507 458
rect 3151 372 3592 373
rect 2818 354 3057 369
rect 3546 357 3592 372
rect 3176 280 3410 326
rect 3456 280 3467 326
rect 3176 279 3467 280
rect 3546 311 3880 357
rect 4302 311 4321 357
rect 2254 215 2432 226
rect 2300 169 2432 215
rect 2511 198 2522 244
rect 2568 198 2842 244
rect 2888 198 2899 244
rect 2254 158 2432 169
rect 1622 106 2208 152
rect 2386 152 2432 158
rect 3176 152 3222 279
rect 3546 167 3592 311
rect 4402 263 4507 412
rect 4009 217 4507 263
rect 2386 106 3222 152
rect 3311 121 3322 167
rect 3368 121 3379 167
rect 3311 60 3379 121
rect 3546 110 3592 121
rect 3770 167 3816 178
rect 3770 60 3816 121
rect 4009 167 4056 217
rect 4402 167 4507 217
rect 4009 121 4010 167
rect 4009 110 4056 121
rect 4223 121 4234 167
rect 4280 121 4291 167
rect 4223 60 4291 121
rect 4402 121 4458 167
rect 4504 121 4507 167
rect 4402 110 4507 121
rect 4682 167 4728 178
rect 4682 60 4728 121
rect 0 -60 4816 60
<< labels >>
flabel metal1 s 578 354 806 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 4334 458 4507 676 0 FreeSans 600 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2818 354 3057 430 0 FreeSans 600 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 724 4816 844 0 FreeSans 600 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1491 210 1559 215 0 FreeSans 600 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 56 353 318 426 0 FreeSans 600 0 0 0 CLK
port 3 nsew clock input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 4010 458 4056 676 1 Q
port 4 nsew default output
rlabel metal1 s 4010 412 4507 458 1 Q
port 4 nsew default output
rlabel metal1 s 4402 263 4507 412 1 Q
port 4 nsew default output
rlabel metal1 s 4009 217 4507 263 1 Q
port 4 nsew default output
rlabel metal1 s 4402 110 4507 217 1 Q
port 4 nsew default output
rlabel metal1 s 4009 110 4056 217 1 Q
port 4 nsew default output
rlabel metal1 s 4682 689 4728 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4234 689 4280 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3750 689 3796 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3341 689 3387 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2859 689 2927 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2055 689 2123 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1535 689 1603 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 689 716 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 689 330 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4682 601 4728 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4234 601 4280 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3750 601 3796 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3341 601 3387 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2859 601 2927 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2055 601 2123 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 601 716 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 601 330 689 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4682 586 4728 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4234 586 4280 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3750 586 3796 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3341 586 3387 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 586 716 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 586 330 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4682 569 4728 586 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4234 569 4280 586 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3750 569 3796 586 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3341 569 3387 586 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 569 716 586 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4682 506 4728 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4234 506 4280 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3750 506 3796 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3341 506 3387 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 630 210 698 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 178 1559 210 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 630 178 698 210 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 178 330 210 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4682 167 4728 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3770 167 3816 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 167 1559 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 630 167 698 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 167 330 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4682 60 4728 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4223 60 4291 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3770 60 3816 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3311 60 3379 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 60 1559 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 630 60 698 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 167 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4816 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 784
string GDS_END 1077356
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1067288
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
