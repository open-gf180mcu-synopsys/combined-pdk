magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1020 1270
<< nmos >>
rect 190 210 250 380
rect 530 210 590 380
rect 730 210 790 380
<< pmos >>
rect 190 720 250 1060
rect 530 720 590 1060
rect 730 720 790 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 430 318 530 380
rect 430 272 452 318
rect 498 272 530 318
rect 430 210 530 272
rect 590 318 730 380
rect 590 272 622 318
rect 668 272 730 318
rect 590 210 730 272
rect 790 318 920 380
rect 790 272 852 318
rect 898 272 920 318
rect 790 210 920 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 350 1060
rect 250 773 282 1007
rect 328 773 350 1007
rect 250 720 350 773
rect 430 1007 530 1060
rect 430 773 452 1007
rect 498 773 530 1007
rect 430 720 530 773
rect 590 1028 730 1060
rect 590 982 622 1028
rect 668 982 730 1028
rect 590 720 730 982
rect 790 1007 920 1060
rect 790 773 852 1007
rect 898 773 920 1007
rect 790 720 920 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 852 272 898 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 452 773 498 1007
rect 622 982 668 1028
rect 852 773 898 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 290 1198 440 1220
rect 290 1152 352 1198
rect 398 1152 440 1198
rect 290 1130 440 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 530 1060 590 1110
rect 730 1060 790 1110
rect 190 670 250 720
rect 120 638 250 670
rect 120 592 142 638
rect 188 600 250 638
rect 530 600 590 720
rect 730 700 790 720
rect 710 678 810 700
rect 710 632 737 678
rect 783 632 810 678
rect 710 610 810 632
rect 188 592 660 600
rect 120 570 660 592
rect 190 560 660 570
rect 190 550 790 560
rect 190 380 250 550
rect 610 510 790 550
rect 300 473 400 500
rect 300 427 327 473
rect 373 460 400 473
rect 373 427 590 460
rect 300 410 590 427
rect 300 400 400 410
rect 530 380 590 410
rect 730 380 790 510
rect 190 160 250 210
rect 530 160 590 210
rect 730 160 790 210
<< polycontact >>
rect 142 592 188 638
rect 737 632 783 678
rect 327 427 373 473
<< metal1 >>
rect 0 1198 1020 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1020 1198
rect 0 1130 1020 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 690 330 773
rect 450 1007 500 1060
rect 450 773 452 1007
rect 498 773 500 1007
rect 280 686 390 690
rect 110 646 210 650
rect 110 594 134 646
rect 186 638 210 646
rect 110 592 142 594
rect 188 592 210 638
rect 110 590 210 592
rect 280 634 314 686
rect 366 634 390 686
rect 280 630 390 634
rect 280 480 330 630
rect 450 530 500 773
rect 620 1028 670 1060
rect 620 982 622 1028
rect 668 982 670 1028
rect 620 930 670 982
rect 850 1007 900 1060
rect 620 906 680 930
rect 620 854 624 906
rect 676 854 680 906
rect 620 830 680 854
rect 450 516 570 530
rect 280 473 400 480
rect 280 427 327 473
rect 373 427 400 473
rect 280 420 400 427
rect 450 464 494 516
rect 546 464 570 516
rect 450 450 570 464
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 420
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 450 318 500 450
rect 450 272 452 318
rect 498 272 500 318
rect 450 210 500 272
rect 620 318 670 830
rect 850 773 852 1007
rect 898 773 900 1007
rect 730 686 790 710
rect 730 634 734 686
rect 786 634 790 686
rect 730 632 737 634
rect 783 632 790 634
rect 730 600 790 632
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 850 530 900 773
rect 850 516 950 530
rect 850 464 874 516
rect 926 464 950 516
rect 850 450 950 464
rect 850 318 900 450
rect 850 272 852 318
rect 898 272 900 318
rect 850 210 900 272
rect 0 118 1020 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1020 118
rect 0 0 1020 72
<< via1 >>
rect 134 638 186 646
rect 134 594 142 638
rect 142 594 186 638
rect 314 634 366 686
rect 624 854 676 906
rect 494 464 546 516
rect 734 678 786 686
rect 734 634 737 678
rect 737 634 783 678
rect 783 634 786 678
rect 874 464 926 516
<< metal2 >>
rect 600 906 700 920
rect 600 854 624 906
rect 676 854 700 906
rect 600 840 700 854
rect 290 690 390 700
rect 710 690 810 700
rect 290 686 810 690
rect 110 646 210 660
rect 110 594 134 646
rect 186 594 210 646
rect 290 634 314 686
rect 366 634 734 686
rect 786 634 810 686
rect 290 630 810 634
rect 290 620 390 630
rect 710 620 810 630
rect 110 580 210 594
rect 470 516 570 530
rect 470 464 494 516
rect 546 464 570 516
rect 470 450 570 464
rect 850 516 950 530
rect 850 464 874 516
rect 926 464 950 516
rect 850 450 950 464
<< labels >>
rlabel via1 s 494 464 546 516 4 A
port 1 nsew signal input
rlabel via1 s 874 464 926 516 4 B
port 2 nsew signal input
rlabel via1 s 134 594 186 646 4 Sel
port 3 nsew signal output
rlabel via1 s 624 854 676 906 4 Y
port 4 nsew signal output
rlabel metal1 s 110 720 160 1270 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 1130 1020 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 0 1020 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 470 450 570 530 1 A
port 1 nsew signal input
rlabel metal1 s 450 210 500 1060 1 A
port 1 nsew signal input
rlabel metal1 s 450 450 570 530 1 A
port 1 nsew signal input
rlabel metal2 s 850 450 950 530 1 B
port 2 nsew signal input
rlabel metal1 s 850 210 900 1060 1 B
port 2 nsew signal input
rlabel metal1 s 850 450 950 530 1 B
port 2 nsew signal input
rlabel metal2 s 110 580 210 660 1 Sel
port 3 nsew signal output
rlabel metal1 s 110 590 210 650 1 Sel
port 3 nsew signal output
rlabel metal2 s 600 840 700 920 1 Y
port 4 nsew signal output
rlabel metal1 s 620 210 670 1060 1 Y
port 4 nsew signal output
rlabel metal1 s 620 830 680 930 1 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1020 1270
string GDS_END 328530
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 321316
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
