magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use npn_00p54x02p00_0  npn_00p54x02p00_0_0
timestamp 1750858719
transform 1 0 1320 0 1 1320
box -1264 -1264 1372 1664
<< labels >>
flabel metal1 s 1325 1325 1325 1325 0 FreeSans 200 0 0 0 I1_default_E
port 3 nsew
flabel metal1 s 61 61 61 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 61 61 61 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 2113 61 2113 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 2613 61 2613 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 61 2905 61 2905 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 1029 1029 1029 1029 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 1645 1029 1645 1029 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 1029 1937 1029 1937 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 1177 1177 1177 1177 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 1497 1177 1497 1177 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 1177 1789 1177 1789 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
<< properties >>
string GDS_END 12842
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_00p54x02p00.gds
string GDS_START 11932
string device primitive
<< end >>
