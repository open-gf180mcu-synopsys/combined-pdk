magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 760 1070 830
rect 145 635 170 760
rect 485 555 510 760
rect 185 453 235 455
rect 185 427 197 453
rect 223 427 235 453
rect 185 425 235 427
rect 740 555 765 760
rect 900 555 925 760
rect 985 525 1010 725
rect 985 520 1025 525
rect 985 518 1035 520
rect 145 70 185 190
rect 470 70 510 190
rect 705 293 755 295
rect 705 267 717 293
rect 743 267 755 293
rect 705 265 755 267
rect 985 492 997 518
rect 1023 492 1035 518
rect 985 490 1035 492
rect 985 485 1025 490
rect 740 70 765 190
rect 900 70 925 190
rect 985 105 1010 485
rect 0 0 1070 70
<< via1 >>
rect 197 427 223 453
rect 717 267 743 293
rect 997 492 1023 518
<< obsm1 >>
rect 60 395 85 725
rect 315 580 340 725
rect 115 555 340 580
rect 570 560 595 725
rect 115 455 140 555
rect 570 535 620 560
rect 260 480 310 510
rect 110 425 155 455
rect 50 390 85 395
rect 35 360 85 390
rect 45 355 85 360
rect 60 105 85 355
rect 115 240 140 425
rect 270 295 300 480
rect 345 425 395 455
rect 520 425 570 455
rect 450 360 500 390
rect 595 295 620 535
rect 655 460 680 725
rect 815 540 840 725
rect 815 520 855 540
rect 815 515 865 520
rect 815 490 950 515
rect 815 485 855 490
rect 655 455 695 460
rect 645 425 695 455
rect 270 265 620 295
rect 115 215 340 240
rect 595 230 620 265
rect 315 105 340 215
rect 570 205 620 230
rect 655 420 695 425
rect 570 105 595 205
rect 655 105 680 420
rect 845 360 895 390
rect 920 240 950 490
rect 815 215 950 240
rect 815 105 840 215
<< metal2 >>
rect 990 520 1030 525
rect 985 518 1035 520
rect 985 492 997 518
rect 1023 492 1035 518
rect 985 490 1035 492
rect 990 485 1030 490
rect 185 453 235 460
rect 185 427 197 453
rect 223 427 235 453
rect 185 420 235 427
rect 705 293 755 300
rect 705 267 717 293
rect 743 267 755 293
rect 705 260 755 267
<< obsm2 >>
rect 820 520 860 525
rect 815 490 865 520
rect 820 485 860 490
rect 350 455 390 460
rect 520 455 570 460
rect 645 455 695 460
rect 345 425 695 455
rect 350 420 390 425
rect 520 420 570 425
rect 645 420 695 425
rect 35 390 85 395
rect 455 390 495 395
rect 845 390 895 395
rect 35 360 895 390
rect 35 355 85 360
rect 455 355 495 360
rect 845 355 895 360
<< labels >>
rlabel metal1 s 145 635 170 830 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 485 555 510 830 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 740 555 765 830 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 900 555 925 830 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 760 1070 830 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 145 0 185 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 470 0 510 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 740 0 765 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 900 0 925 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1070 70 6 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 717 267 743 293 6 CLK
port 3 nsew clock input
rlabel metal2 s 705 260 755 300 6 CLK
port 3 nsew clock input
rlabel metal1 s 705 265 755 295 6 CLK
port 3 nsew clock input
rlabel via1 s 197 427 223 453 6 D
port 1 nsew signal input
rlabel metal2 s 185 420 235 460 6 D
port 1 nsew signal input
rlabel metal1 s 185 425 235 455 6 D
port 1 nsew signal input
rlabel via1 s 997 492 1023 518 6 Q
port 2 nsew signal output
rlabel metal2 s 990 485 1030 525 6 Q
port 2 nsew signal output
rlabel metal2 s 985 490 1035 520 6 Q
port 2 nsew signal output
rlabel metal1 s 985 105 1010 725 6 Q
port 2 nsew signal output
rlabel metal1 s 985 485 1025 525 6 Q
port 2 nsew signal output
rlabel metal1 s 985 490 1035 520 6 Q
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1070 830
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 403594
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 388226
<< end >>
