VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__fill5
  CLASS PAD SPACER ;
  FOREIGN gf180mcu_fd_io__fill5 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 1.730 134.000 5.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 150.000 5.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 166.000 5.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 182.000 5.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 214.000 5.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 118.000 5.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 206.000 5.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 262.000 5.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 270.000 5.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 278.000 5.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 294.000 5.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 1.730 334.000 5.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 1.450 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 1.450 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 1.450 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 1.450 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 1.450 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 1.450 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 1.450 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 1.450 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 1.450 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 1.450 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 1.450 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 1.450 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 3.610 70.000 5.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 86.000 5.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 102.000 5.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 230.000 5.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 126.000 5.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 198.000 5.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 286.000 5.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 302.000 5.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 326.000 5.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 3.610 342.000 5.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 3.330 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 3.330 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 3.330 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 3.330 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 3.330 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 3.330 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 3.330 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 3.330 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 3.330 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 3.330 85.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 2.690 254.000 5.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 2.690 310.000 5.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 2.410 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 2.410 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 4.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 4.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 5.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 67.350 5.000 348.300 ;
  END
END gf180mcu_fd_io__fill5
END LIBRARY

