magic
tech gf180mcuA
timestamp 1750858719
<< properties >>
string FIXED_BBOX 0 0 8 166
string GDS_END 404614
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 404338
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
