magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 2260 1270
<< nmos >>
rect 200 210 260 380
rect 400 210 460 380
rect 540 210 600 380
rect 710 210 770 380
rect 950 210 1010 380
rect 1150 210 1210 380
rect 1510 210 1570 380
rect 1830 210 1890 380
rect 2000 210 2060 380
<< pmos >>
rect 200 720 260 1060
rect 370 720 430 1060
rect 540 720 600 1060
rect 710 720 770 1060
rect 980 720 1040 1060
rect 1150 720 1210 1060
rect 1510 720 1570 1060
rect 1830 720 1890 1060
rect 2000 720 2060 1060
<< ndiff >>
rect 100 318 200 380
rect 100 272 122 318
rect 168 272 200 318
rect 100 210 200 272
rect 260 288 400 380
rect 260 242 307 288
rect 353 242 400 288
rect 260 210 400 242
rect 460 210 540 380
rect 600 293 710 380
rect 600 247 632 293
rect 678 247 710 293
rect 600 210 710 247
rect 770 210 950 380
rect 1010 283 1150 380
rect 1010 237 1057 283
rect 1103 237 1150 283
rect 1010 210 1150 237
rect 1210 318 1310 380
rect 1210 272 1242 318
rect 1288 272 1310 318
rect 1210 210 1310 272
rect 1410 318 1510 380
rect 1410 272 1432 318
rect 1478 272 1510 318
rect 1410 210 1510 272
rect 1570 318 1670 380
rect 1570 272 1602 318
rect 1648 272 1670 318
rect 1570 210 1670 272
rect 1730 318 1830 380
rect 1730 272 1752 318
rect 1798 272 1830 318
rect 1730 210 1830 272
rect 1890 283 2000 380
rect 1890 237 1922 283
rect 1968 237 2000 283
rect 1890 210 2000 237
rect 2060 318 2160 380
rect 2060 272 2092 318
rect 2138 272 2160 318
rect 2060 210 2160 272
<< pdiff >>
rect 100 1007 200 1060
rect 100 773 122 1007
rect 168 773 200 1007
rect 100 720 200 773
rect 260 1040 370 1060
rect 260 900 292 1040
rect 338 900 370 1040
rect 260 720 370 900
rect 430 720 540 1060
rect 600 1037 710 1060
rect 600 803 632 1037
rect 678 803 710 1037
rect 600 720 710 803
rect 770 720 980 1060
rect 1040 1032 1150 1060
rect 1040 798 1072 1032
rect 1118 798 1150 1032
rect 1040 720 1150 798
rect 1210 1037 1310 1060
rect 1210 803 1242 1037
rect 1288 803 1310 1037
rect 1210 720 1310 803
rect 1410 1005 1510 1060
rect 1410 865 1432 1005
rect 1478 865 1510 1005
rect 1410 720 1510 865
rect 1570 1012 1670 1060
rect 1570 778 1602 1012
rect 1648 778 1670 1012
rect 1570 720 1670 778
rect 1730 1012 1830 1060
rect 1730 778 1752 1012
rect 1798 778 1830 1012
rect 1730 720 1830 778
rect 1890 1030 2000 1060
rect 1890 890 1922 1030
rect 1968 890 2000 1030
rect 1890 720 2000 890
rect 2060 1007 2160 1060
rect 2060 773 2092 1007
rect 2138 773 2160 1007
rect 2060 720 2160 773
<< ndiffc >>
rect 122 272 168 318
rect 307 242 353 288
rect 632 247 678 293
rect 1057 237 1103 283
rect 1242 272 1288 318
rect 1432 272 1478 318
rect 1602 272 1648 318
rect 1752 272 1798 318
rect 1922 237 1968 283
rect 2092 272 2138 318
<< pdiffc >>
rect 122 773 168 1007
rect 292 900 338 1040
rect 632 803 678 1037
rect 1072 798 1118 1032
rect 1242 803 1288 1037
rect 1432 865 1478 1005
rect 1602 778 1648 1012
rect 1752 778 1798 1012
rect 1922 890 1968 1030
rect 2092 773 2138 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1030 118 1180 140
rect 1030 72 1082 118
rect 1128 72 1180 118
rect 1030 50 1180 72
rect 1280 118 1430 140
rect 1280 72 1332 118
rect 1378 72 1430 118
rect 1280 50 1430 72
rect 1530 118 1680 140
rect 1530 72 1582 118
rect 1628 72 1680 118
rect 1530 50 1680 72
rect 1780 118 1930 140
rect 1780 72 1832 118
rect 1878 72 1930 118
rect 1780 50 1930 72
rect 2030 118 2180 140
rect 2030 72 2082 118
rect 2128 72 2180 118
rect 2030 50 2180 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 310 1198 460 1220
rect 310 1152 362 1198
rect 408 1152 460 1198
rect 310 1130 460 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1030 1198 1180 1220
rect 1030 1152 1082 1198
rect 1128 1152 1180 1198
rect 1030 1130 1180 1152
rect 1280 1198 1430 1220
rect 1280 1152 1332 1198
rect 1378 1152 1430 1198
rect 1280 1130 1430 1152
rect 1530 1198 1680 1220
rect 1530 1152 1582 1198
rect 1628 1152 1680 1198
rect 1530 1130 1680 1152
rect 1780 1198 1930 1220
rect 1780 1152 1832 1198
rect 1878 1152 1930 1198
rect 1780 1130 1930 1152
rect 2030 1198 2180 1220
rect 2030 1152 2082 1198
rect 2128 1152 2180 1198
rect 2030 1130 2180 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 592 72 638 118
rect 832 72 878 118
rect 1082 72 1128 118
rect 1332 72 1378 118
rect 1582 72 1628 118
rect 1832 72 1878 118
rect 2082 72 2128 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 362 1152 408 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1082 1152 1128 1198
rect 1332 1152 1378 1198
rect 1582 1152 1628 1198
rect 1832 1152 1878 1198
rect 2082 1152 2128 1198
<< polysilicon >>
rect 200 1060 260 1110
rect 370 1060 430 1110
rect 540 1060 600 1110
rect 710 1060 770 1110
rect 980 1060 1040 1110
rect 1150 1060 1210 1110
rect 1510 1060 1570 1110
rect 1830 1060 1890 1110
rect 2000 1060 2060 1110
rect 200 700 260 720
rect 200 673 320 700
rect 200 627 237 673
rect 283 627 320 673
rect 200 600 320 627
rect 370 670 430 720
rect 540 700 600 720
rect 710 700 770 720
rect 520 673 620 700
rect 370 643 470 670
rect 200 380 260 600
rect 370 597 397 643
rect 443 597 470 643
rect 520 627 547 673
rect 593 627 620 673
rect 520 600 620 627
rect 680 673 780 700
rect 680 627 707 673
rect 753 627 780 673
rect 680 600 780 627
rect 370 570 470 597
rect 370 440 430 570
rect 710 550 770 600
rect 540 510 770 550
rect 830 563 930 590
rect 830 517 857 563
rect 903 517 930 563
rect 370 400 460 440
rect 400 380 460 400
rect 540 380 600 510
rect 830 490 930 517
rect 980 570 1040 720
rect 1150 700 1210 720
rect 1140 673 1240 700
rect 1140 627 1167 673
rect 1213 627 1240 673
rect 1140 600 1240 627
rect 1510 670 1570 720
rect 1510 648 1640 670
rect 1510 602 1572 648
rect 1618 602 1640 648
rect 980 543 1100 570
rect 980 497 1027 543
rect 1073 497 1100 543
rect 830 460 900 490
rect 710 420 900 460
rect 980 470 1100 497
rect 980 440 1040 470
rect 710 380 770 420
rect 950 400 1040 440
rect 950 380 1010 400
rect 1150 380 1210 600
rect 1510 580 1640 602
rect 1510 380 1570 580
rect 1830 570 1890 720
rect 2000 570 2060 720
rect 1800 548 1890 570
rect 1800 502 1822 548
rect 1868 502 1890 548
rect 1800 480 1890 502
rect 1830 380 1890 480
rect 1940 543 2060 570
rect 1940 497 1967 543
rect 2013 497 2060 543
rect 1940 470 2060 497
rect 2000 380 2060 470
rect 200 160 260 210
rect 400 160 460 210
rect 540 160 600 210
rect 710 160 770 210
rect 950 160 1010 210
rect 1150 160 1210 210
rect 1510 160 1570 210
rect 1830 160 1890 210
rect 2000 160 2060 210
<< polycontact >>
rect 237 627 283 673
rect 397 597 443 643
rect 547 627 593 673
rect 707 627 753 673
rect 857 517 903 563
rect 1167 627 1213 673
rect 1572 602 1618 648
rect 1027 497 1073 543
rect 1822 502 1868 548
rect 1967 497 2013 543
<< metal1 >>
rect 0 1198 2260 1270
rect 0 1152 112 1198
rect 158 1152 362 1198
rect 408 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1082 1198
rect 1128 1152 1332 1198
rect 1378 1152 1582 1198
rect 1628 1152 1832 1198
rect 1878 1152 2082 1198
rect 2128 1152 2260 1198
rect 0 1130 2260 1152
rect 120 1007 170 1060
rect 120 773 122 1007
rect 168 773 170 1007
rect 290 1040 340 1130
rect 290 900 292 1040
rect 338 900 340 1040
rect 290 880 340 900
rect 630 1037 680 1060
rect 630 830 632 1037
rect 120 530 170 773
rect 230 803 632 830
rect 678 803 680 1037
rect 230 780 680 803
rect 1070 1032 1120 1130
rect 1070 798 1072 1032
rect 1118 798 1120 1032
rect 230 680 280 780
rect 1070 770 1120 798
rect 1240 1037 1290 1060
rect 1240 803 1242 1037
rect 1288 803 1290 1037
rect 1240 800 1290 803
rect 1430 1005 1480 1060
rect 1430 865 1432 1005
rect 1478 865 1480 1005
rect 1240 750 1340 800
rect 220 673 310 680
rect 220 627 237 673
rect 283 627 310 673
rect 520 673 620 680
rect 220 620 310 627
rect 370 646 470 650
rect 100 520 170 530
rect 70 516 170 520
rect 70 464 94 516
rect 146 464 170 516
rect 70 460 170 464
rect 90 450 170 460
rect 120 318 170 450
rect 230 450 280 620
rect 370 594 394 646
rect 446 594 470 646
rect 520 627 547 673
rect 593 627 620 673
rect 520 620 620 627
rect 680 673 780 680
rect 680 646 707 673
rect 753 646 780 673
rect 370 590 470 594
rect 540 540 600 620
rect 680 594 704 646
rect 756 594 780 646
rect 1140 676 1240 680
rect 1140 624 1164 676
rect 1216 624 1240 676
rect 1140 620 1240 624
rect 680 590 780 594
rect 830 563 930 570
rect 830 540 857 563
rect 540 517 857 540
rect 903 517 930 563
rect 540 510 930 517
rect 1000 546 1100 550
rect 540 490 910 510
rect 1000 494 1024 546
rect 1076 494 1100 546
rect 1000 490 1100 494
rect 540 480 900 490
rect 230 400 480 450
rect 120 272 122 318
rect 168 272 170 318
rect 120 210 170 272
rect 290 288 370 320
rect 290 242 307 288
rect 353 242 370 288
rect 430 310 480 400
rect 840 410 900 480
rect 1290 470 1340 750
rect 1430 680 1480 865
rect 1600 1012 1650 1130
rect 1600 778 1602 1012
rect 1648 778 1650 1012
rect 1600 730 1650 778
rect 1750 1012 1800 1060
rect 1750 778 1752 1012
rect 1798 778 1800 1012
rect 1920 1030 1970 1130
rect 1920 890 1922 1030
rect 1968 890 1970 1030
rect 1920 860 1970 890
rect 2090 1007 2140 1060
rect 1750 740 1800 778
rect 2090 773 2092 1007
rect 2138 773 2140 1007
rect 1750 690 2020 740
rect 1390 676 1490 680
rect 1390 624 1414 676
rect 1466 624 1490 676
rect 1390 620 1490 624
rect 1550 648 1650 650
rect 1240 420 1340 470
rect 1240 410 1290 420
rect 840 360 1290 410
rect 630 310 680 330
rect 1240 318 1290 360
rect 430 293 680 310
rect 430 260 632 293
rect 290 140 370 242
rect 630 247 632 260
rect 678 247 680 293
rect 630 210 680 247
rect 1040 283 1120 310
rect 1040 237 1057 283
rect 1103 237 1120 283
rect 1040 140 1120 237
rect 1240 272 1242 318
rect 1288 272 1290 318
rect 1240 210 1290 272
rect 1430 318 1480 620
rect 1550 602 1572 648
rect 1618 646 1650 648
rect 1550 594 1574 602
rect 1626 594 1650 646
rect 1550 590 1650 594
rect 1800 548 1900 550
rect 1800 502 1822 548
rect 1868 546 1900 548
rect 1800 494 1824 502
rect 1876 494 1900 546
rect 1800 490 1900 494
rect 1960 543 2020 690
rect 1960 497 1967 543
rect 2013 497 2020 543
rect 1960 440 2020 497
rect 1750 390 2020 440
rect 2090 660 2140 773
rect 2090 650 2170 660
rect 2090 646 2190 650
rect 2090 594 2114 646
rect 2166 594 2190 646
rect 2090 590 2190 594
rect 2090 580 2170 590
rect 1430 272 1432 318
rect 1478 272 1480 318
rect 1430 210 1480 272
rect 1600 318 1650 380
rect 1600 272 1602 318
rect 1648 272 1650 318
rect 1600 140 1650 272
rect 1750 318 1800 390
rect 1750 272 1752 318
rect 1798 272 1800 318
rect 2090 318 2140 580
rect 1750 210 1800 272
rect 1920 283 1970 310
rect 1920 237 1922 283
rect 1968 237 1970 283
rect 1920 140 1970 237
rect 2090 272 2092 318
rect 2138 272 2140 318
rect 2090 210 2140 272
rect 0 118 2260 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 592 118
rect 638 72 832 118
rect 878 72 1082 118
rect 1128 72 1332 118
rect 1378 72 1582 118
rect 1628 72 1832 118
rect 1878 72 2082 118
rect 2128 72 2260 118
rect 0 0 2260 72
<< via1 >>
rect 94 464 146 516
rect 394 643 446 646
rect 394 597 397 643
rect 397 597 443 643
rect 443 597 446 643
rect 394 594 446 597
rect 704 627 707 646
rect 707 627 753 646
rect 753 627 756 646
rect 704 594 756 627
rect 1164 673 1216 676
rect 1164 627 1167 673
rect 1167 627 1213 673
rect 1213 627 1216 673
rect 1164 624 1216 627
rect 1024 543 1076 546
rect 1024 497 1027 543
rect 1027 497 1073 543
rect 1073 497 1076 543
rect 1024 494 1076 497
rect 1414 624 1466 676
rect 1574 602 1618 646
rect 1618 602 1626 646
rect 1574 594 1626 602
rect 1824 502 1868 546
rect 1868 502 1876 546
rect 1824 494 1876 502
rect 2114 594 2166 646
<< metal2 >>
rect 1140 680 1240 690
rect 1390 680 1490 690
rect 700 676 1490 680
rect 700 660 1164 676
rect 370 646 470 660
rect 690 650 1164 660
rect 370 594 394 646
rect 446 594 470 646
rect 370 580 470 594
rect 680 646 1164 650
rect 680 594 704 646
rect 756 624 1164 646
rect 1216 624 1414 676
rect 1466 624 1490 676
rect 756 620 1490 624
rect 756 594 780 620
rect 1140 610 1240 620
rect 1390 610 1490 620
rect 1550 646 1650 660
rect 2100 650 2180 660
rect 680 590 780 594
rect 1550 594 1574 646
rect 1626 594 1650 646
rect 690 580 770 590
rect 1550 580 1650 594
rect 2090 646 2190 650
rect 2090 594 2114 646
rect 2166 594 2190 646
rect 2090 590 2190 594
rect 2100 580 2180 590
rect 1010 550 1100 560
rect 1800 550 1900 560
rect 920 546 1100 550
rect 70 520 170 530
rect 920 520 1024 546
rect 70 516 1024 520
rect 70 464 94 516
rect 146 494 1024 516
rect 1076 510 1100 546
rect 1790 546 1900 550
rect 1790 510 1824 546
rect 1076 494 1824 510
rect 1876 494 1900 546
rect 146 480 1900 494
rect 146 464 980 480
rect 70 460 980 464
rect 70 450 170 460
rect 1040 450 1850 480
<< labels >>
rlabel via1 s 394 594 446 646 4 D
port 1 nsew signal input
rlabel via1 s 2114 594 2166 646 4 Q
port 2 nsew signal output
rlabel via1 s 1574 594 1626 646 4 CLK
port 3 nsew clock input
rlabel metal1 s 290 880 340 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 0 370 320 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1070 770 1120 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1600 730 1650 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1920 860 1970 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 2260 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1040 0 1120 310 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1600 0 1650 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1920 0 1970 310 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2260 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 1550 580 1650 660 1 CLK
port 3 nsew clock input
rlabel metal1 s 1550 590 1650 650 1 CLK
port 3 nsew clock input
rlabel metal2 s 370 580 470 660 1 D
port 1 nsew signal input
rlabel metal1 s 370 590 470 650 1 D
port 1 nsew signal input
rlabel metal2 s 2100 580 2180 660 1 Q
port 2 nsew signal output
rlabel metal2 s 2090 590 2190 650 1 Q
port 2 nsew signal output
rlabel metal1 s 2090 210 2140 1060 1 Q
port 2 nsew signal output
rlabel metal1 s 2090 580 2170 660 1 Q
port 2 nsew signal output
rlabel metal1 s 2090 590 2190 650 1 Q
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2260 1270
string GDS_END 282408
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 266080
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
