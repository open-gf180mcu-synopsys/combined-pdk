magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 377 4006 870
rect -86 352 2018 377
rect 3590 352 4006 377
<< pwell >>
rect -86 -86 4006 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2184 93 2304 257
rect 2408 93 2528 257
rect 2632 93 2752 257
rect 2856 93 2976 257
rect 3080 93 3200 257
rect 3304 93 3424 257
rect 3572 68 3692 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 572 497 672 716
rect 816 497 916 716
rect 1020 497 1120 716
rect 1264 497 1364 716
rect 1468 497 1568 716
rect 1692 497 1792 716
rect 1936 497 2036 716
rect 2204 497 2304 716
rect 2408 497 2508 716
rect 2652 497 2752 716
rect 2856 497 2956 716
rect 3100 497 3200 716
rect 3304 497 3404 716
rect 3572 497 3672 716
<< mvndiff >>
rect 2096 244 2184 257
rect 2096 232 2109 244
rect 36 156 124 232
rect 36 110 49 156
rect 95 110 124 156
rect 36 68 124 110
rect 244 143 348 232
rect 244 97 273 143
rect 319 97 348 143
rect 244 68 348 97
rect 468 156 572 232
rect 468 110 497 156
rect 543 110 572 156
rect 468 68 572 110
rect 692 143 796 232
rect 692 97 721 143
rect 767 97 796 143
rect 692 68 796 97
rect 916 156 1020 232
rect 916 110 945 156
rect 991 110 1020 156
rect 916 68 1020 110
rect 1140 143 1244 232
rect 1140 97 1169 143
rect 1215 97 1244 143
rect 1140 68 1244 97
rect 1364 156 1468 232
rect 1364 110 1393 156
rect 1439 110 1468 156
rect 1364 68 1468 110
rect 1588 143 1692 232
rect 1588 97 1617 143
rect 1663 97 1692 143
rect 1588 68 1692 97
rect 1812 152 1916 232
rect 1812 106 1841 152
rect 1887 106 1916 152
rect 1812 68 1916 106
rect 2036 198 2109 232
rect 2155 198 2184 244
rect 2036 93 2184 198
rect 2304 152 2408 257
rect 2304 106 2333 152
rect 2379 106 2408 152
rect 2304 93 2408 106
rect 2528 244 2632 257
rect 2528 198 2557 244
rect 2603 198 2632 244
rect 2528 93 2632 198
rect 2752 152 2856 257
rect 2752 106 2781 152
rect 2827 106 2856 152
rect 2752 93 2856 106
rect 2976 244 3080 257
rect 2976 198 3005 244
rect 3051 198 3080 244
rect 2976 93 3080 198
rect 3200 152 3304 257
rect 3200 106 3229 152
rect 3275 106 3304 152
rect 3200 93 3304 106
rect 3424 244 3512 257
rect 3424 198 3453 244
rect 3499 232 3512 244
rect 3499 198 3572 232
rect 3424 93 3572 198
rect 2036 68 2116 93
rect 3492 68 3572 93
rect 3692 152 3780 232
rect 3692 106 3721 152
rect 3767 106 3780 152
rect 3692 68 3780 106
<< mvpdiff >>
rect 56 677 144 716
rect 56 537 69 677
rect 115 537 144 677
rect 56 497 144 537
rect 244 497 368 716
rect 468 639 572 716
rect 468 593 497 639
rect 543 593 572 639
rect 468 497 572 593
rect 672 497 816 716
rect 916 697 1020 716
rect 916 651 945 697
rect 991 651 1020 697
rect 916 497 1020 651
rect 1120 497 1264 716
rect 1364 665 1468 716
rect 1364 525 1393 665
rect 1439 525 1468 665
rect 1364 497 1468 525
rect 1568 497 1692 716
rect 1792 697 1936 716
rect 1792 651 1841 697
rect 1887 651 1936 697
rect 1792 497 1936 651
rect 2036 497 2204 716
rect 2304 639 2408 716
rect 2304 593 2333 639
rect 2379 593 2408 639
rect 2304 497 2408 593
rect 2508 497 2652 716
rect 2752 697 2856 716
rect 2752 651 2781 697
rect 2827 651 2856 697
rect 2752 497 2856 651
rect 2956 497 3100 716
rect 3200 665 3304 716
rect 3200 525 3229 665
rect 3275 525 3304 665
rect 3200 497 3304 525
rect 3404 497 3572 716
rect 3672 677 3760 716
rect 3672 537 3701 677
rect 3747 537 3760 677
rect 3672 497 3760 537
<< mvndiffc >>
rect 49 110 95 156
rect 273 97 319 143
rect 497 110 543 156
rect 721 97 767 143
rect 945 110 991 156
rect 1169 97 1215 143
rect 1393 110 1439 156
rect 1617 97 1663 143
rect 1841 106 1887 152
rect 2109 198 2155 244
rect 2333 106 2379 152
rect 2557 198 2603 244
rect 2781 106 2827 152
rect 3005 198 3051 244
rect 3229 106 3275 152
rect 3453 198 3499 244
rect 3721 106 3767 152
<< mvpdiffc >>
rect 69 537 115 677
rect 497 593 543 639
rect 945 651 991 697
rect 1393 525 1439 665
rect 1841 651 1887 697
rect 2333 593 2379 639
rect 2781 651 2827 697
rect 3229 525 3275 665
rect 3701 537 3747 677
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 1020 716 1120 760
rect 1264 716 1364 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1936 716 2036 760
rect 2204 716 2304 760
rect 2408 716 2508 760
rect 2652 716 2752 760
rect 2856 716 2956 760
rect 3100 716 3200 760
rect 3304 716 3404 760
rect 3572 716 3672 760
rect 144 401 244 497
rect 368 413 468 497
rect 368 401 395 413
rect 124 382 244 401
rect 124 336 178 382
rect 224 336 244 382
rect 124 232 244 336
rect 348 367 395 401
rect 441 401 468 413
rect 572 413 672 497
rect 572 401 599 413
rect 441 367 599 401
rect 645 401 672 413
rect 816 419 916 497
rect 816 401 843 419
rect 645 367 692 401
rect 348 344 692 367
rect 348 232 468 344
rect 572 232 692 344
rect 796 373 843 401
rect 889 401 916 419
rect 1020 419 1120 497
rect 1020 401 1047 419
rect 889 373 1047 401
rect 1093 401 1120 419
rect 1264 401 1364 497
rect 1468 401 1568 497
rect 1692 419 1792 497
rect 1093 373 1140 401
rect 796 344 1140 373
rect 796 232 916 344
rect 1020 232 1140 344
rect 1244 344 1588 401
rect 1244 327 1364 344
rect 1244 281 1281 327
rect 1327 281 1364 327
rect 1244 232 1364 281
rect 1468 327 1588 344
rect 1468 281 1505 327
rect 1551 281 1588 327
rect 1468 232 1588 281
rect 1692 373 1713 419
rect 1759 401 1792 419
rect 1936 415 2036 497
rect 1936 401 1961 415
rect 1759 373 1812 401
rect 1692 232 1812 373
rect 1916 369 1961 401
rect 2007 369 2036 415
rect 2204 413 2304 497
rect 2204 401 2231 413
rect 1916 232 2036 369
rect 2184 367 2231 401
rect 2277 401 2304 413
rect 2408 413 2508 497
rect 2408 401 2435 413
rect 2277 367 2435 401
rect 2481 401 2508 413
rect 2652 428 2752 497
rect 2652 401 2679 428
rect 2481 367 2528 401
rect 2184 344 2528 367
rect 2184 257 2304 344
rect 2408 257 2528 344
rect 2632 382 2679 401
rect 2725 401 2752 428
rect 2856 428 2956 497
rect 2856 401 2883 428
rect 2725 382 2883 401
rect 2929 401 2956 428
rect 3100 401 3200 497
rect 3304 401 3404 497
rect 3572 428 3672 497
rect 2929 382 2976 401
rect 2632 344 2976 382
rect 2632 257 2752 344
rect 2856 257 2976 344
rect 3080 344 3424 401
rect 3080 336 3200 344
rect 3080 290 3117 336
rect 3163 290 3200 336
rect 3080 257 3200 290
rect 3304 336 3424 344
rect 3304 290 3341 336
rect 3387 290 3424 336
rect 3304 257 3424 290
rect 3572 382 3599 428
rect 3645 401 3672 428
rect 3645 382 3692 401
rect 3572 232 3692 382
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2184 24 2304 93
rect 2408 24 2528 93
rect 2632 24 2752 93
rect 2856 24 2976 93
rect 3080 24 3200 93
rect 3304 24 3424 93
rect 3572 24 3692 68
<< polycontact >>
rect 178 336 224 382
rect 395 367 441 413
rect 599 367 645 413
rect 843 373 889 419
rect 1047 373 1093 419
rect 1281 281 1327 327
rect 1505 281 1551 327
rect 1713 373 1759 419
rect 1961 369 2007 415
rect 2231 367 2277 413
rect 2435 367 2481 413
rect 2679 382 2725 428
rect 2883 382 2929 428
rect 3117 290 3163 336
rect 3341 290 3387 336
rect 3599 382 3645 428
<< metal1 >>
rect 0 724 3920 844
rect 69 677 115 724
rect 934 697 1002 724
rect 934 651 945 697
rect 991 651 1002 697
rect 1830 697 1898 724
rect 1051 665 1781 676
rect 346 639 884 648
rect 346 593 497 639
rect 543 605 884 639
rect 1051 605 1393 665
rect 543 593 1393 605
rect 346 584 1393 593
rect 834 559 1393 584
rect 69 518 115 537
rect 165 472 788 536
rect 1382 525 1393 559
rect 1439 605 1781 665
rect 1830 651 1841 697
rect 1887 651 1898 697
rect 2770 697 2838 724
rect 2770 651 2781 697
rect 2827 651 2838 697
rect 3701 677 3747 724
rect 2888 665 3275 676
rect 1948 639 2721 648
rect 1948 605 2333 639
rect 1439 593 2333 605
rect 2379 605 2721 639
rect 2888 605 3229 665
rect 2379 593 3229 605
rect 1439 584 3229 593
rect 1439 559 1998 584
rect 2671 559 2938 584
rect 1439 525 1450 559
rect 1382 514 1450 525
rect 165 382 229 472
rect 165 336 178 382
rect 224 336 229 382
rect 306 413 672 424
rect 306 367 395 413
rect 441 367 599 413
rect 645 367 672 413
rect 738 419 788 472
rect 738 373 843 419
rect 889 373 1047 419
rect 1093 373 1713 419
rect 1759 373 1770 419
rect 306 357 672 367
rect 165 317 229 336
rect 622 327 672 357
rect 622 281 1281 327
rect 1327 281 1505 327
rect 1551 281 1588 327
rect 1816 244 1876 559
rect 2040 472 2625 536
rect 3229 497 3275 525
rect 3701 518 3747 537
rect 2040 424 2100 472
rect 2575 428 2625 472
rect 1922 415 2100 424
rect 1922 369 1961 415
rect 2007 369 2100 415
rect 1922 360 2100 369
rect 2146 413 2508 424
rect 2146 367 2231 413
rect 2277 367 2435 413
rect 2481 367 2508 413
rect 2575 382 2679 428
rect 2725 382 2883 428
rect 2929 382 3599 428
rect 3645 382 3692 428
rect 2146 357 2508 367
rect 2458 336 2508 357
rect 2458 290 3117 336
rect 3163 290 3341 336
rect 3387 290 3424 336
rect 38 189 1768 235
rect 1816 198 2109 244
rect 2155 198 2557 244
rect 2603 198 3005 244
rect 3051 198 3453 244
rect 3499 198 3512 244
rect 38 156 106 189
rect 38 110 49 156
rect 95 110 106 156
rect 486 156 554 189
rect 262 97 273 143
rect 319 97 330 143
rect 486 110 497 156
rect 543 110 554 156
rect 934 156 1002 189
rect 262 60 330 97
rect 710 97 721 143
rect 767 97 778 143
rect 934 110 945 156
rect 991 110 1002 156
rect 1382 156 1450 189
rect 710 60 778 97
rect 1158 97 1169 143
rect 1215 97 1226 143
rect 1382 110 1393 156
rect 1439 110 1450 156
rect 1722 152 1768 189
rect 1158 60 1226 97
rect 1606 97 1617 143
rect 1663 97 1674 143
rect 1722 106 1841 152
rect 1887 106 2333 152
rect 2379 106 2781 152
rect 2827 106 3229 152
rect 3275 106 3721 152
rect 3767 106 3780 152
rect 1606 60 1674 97
rect 0 -60 3920 60
<< labels >>
flabel metal1 s 306 357 672 424 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 0 724 3920 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1606 60 1674 143 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 2888 648 3275 676 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 2146 357 2508 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 2040 472 2625 536 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel metal1 s 165 472 788 536 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 2458 336 2508 357 1 A1
port 1 nsew default input
rlabel metal1 s 2458 290 3424 336 1 A1
port 1 nsew default input
rlabel metal1 s 2575 428 2625 472 1 A2
port 2 nsew default input
rlabel metal1 s 2040 428 2100 472 1 A2
port 2 nsew default input
rlabel metal1 s 2575 424 3692 428 1 A2
port 2 nsew default input
rlabel metal1 s 2040 424 2100 428 1 A2
port 2 nsew default input
rlabel metal1 s 2575 382 3692 424 1 A2
port 2 nsew default input
rlabel metal1 s 1922 382 2100 424 1 A2
port 2 nsew default input
rlabel metal1 s 1922 360 2100 382 1 A2
port 2 nsew default input
rlabel metal1 s 622 327 672 357 1 B1
port 3 nsew default input
rlabel metal1 s 622 281 1588 327 1 B1
port 3 nsew default input
rlabel metal1 s 738 419 788 472 1 B2
port 4 nsew default input
rlabel metal1 s 165 419 229 472 1 B2
port 4 nsew default input
rlabel metal1 s 738 373 1770 419 1 B2
port 4 nsew default input
rlabel metal1 s 165 373 229 419 1 B2
port 4 nsew default input
rlabel metal1 s 165 317 229 373 1 B2
port 4 nsew default input
rlabel metal1 s 1051 648 1781 676 1 ZN
port 5 nsew default output
rlabel metal1 s 2888 605 3275 648 1 ZN
port 5 nsew default output
rlabel metal1 s 1948 605 2721 648 1 ZN
port 5 nsew default output
rlabel metal1 s 1051 605 1781 648 1 ZN
port 5 nsew default output
rlabel metal1 s 346 605 884 648 1 ZN
port 5 nsew default output
rlabel metal1 s 346 584 3275 605 1 ZN
port 5 nsew default output
rlabel metal1 s 3229 559 3275 584 1 ZN
port 5 nsew default output
rlabel metal1 s 2671 559 2938 584 1 ZN
port 5 nsew default output
rlabel metal1 s 834 559 1998 584 1 ZN
port 5 nsew default output
rlabel metal1 s 3229 514 3275 559 1 ZN
port 5 nsew default output
rlabel metal1 s 1816 514 1876 559 1 ZN
port 5 nsew default output
rlabel metal1 s 1382 514 1450 559 1 ZN
port 5 nsew default output
rlabel metal1 s 3229 497 3275 514 1 ZN
port 5 nsew default output
rlabel metal1 s 1816 497 1876 514 1 ZN
port 5 nsew default output
rlabel metal1 s 1816 244 1876 497 1 ZN
port 5 nsew default output
rlabel metal1 s 1816 198 3512 244 1 ZN
port 5 nsew default output
rlabel metal1 s 3701 651 3747 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2770 651 2838 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1830 651 1898 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 934 651 1002 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 651 115 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3701 518 3747 651 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 518 115 651 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1158 60 1226 143 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 710 60 778 143 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 143 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3920 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 784
string GDS_END 35834
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 28668
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
