magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 800 1270
<< nmos >>
rect 180 210 240 380
rect 350 210 410 380
rect 540 210 600 380
<< pmos >>
rect 210 720 270 1060
rect 330 720 390 1060
rect 520 720 580 1060
<< ndiff >>
rect 80 288 180 380
rect 80 242 102 288
rect 148 242 180 288
rect 80 210 180 242
rect 240 278 350 380
rect 240 232 272 278
rect 318 232 350 278
rect 240 210 350 232
rect 410 288 540 380
rect 410 242 452 288
rect 498 242 540 288
rect 410 210 540 242
rect 600 308 700 380
rect 600 262 632 308
rect 678 262 700 308
rect 600 210 700 262
<< pdiff >>
rect 110 1007 210 1060
rect 110 773 132 1007
rect 178 773 210 1007
rect 110 720 210 773
rect 270 720 330 1060
rect 390 1000 520 1060
rect 390 860 432 1000
rect 478 860 520 1000
rect 390 720 520 860
rect 580 1008 680 1060
rect 580 962 612 1008
rect 658 962 680 1008
rect 580 790 680 962
rect 580 720 690 790
<< ndiffc >>
rect 102 242 148 288
rect 272 232 318 278
rect 452 242 498 288
rect 632 262 678 308
<< pdiffc >>
rect 132 773 178 1007
rect 432 860 478 1000
rect 612 962 658 1008
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
<< polysilicon >>
rect 210 1060 270 1110
rect 330 1060 390 1110
rect 520 1060 580 1110
rect 210 700 270 720
rect 160 660 270 700
rect 330 670 390 720
rect 160 540 220 660
rect 320 643 430 670
rect 320 597 357 643
rect 403 597 430 643
rect 320 570 430 597
rect 110 513 220 540
rect 110 467 147 513
rect 193 470 220 513
rect 330 470 390 570
rect 520 540 580 720
rect 470 513 600 540
rect 193 467 240 470
rect 110 440 240 467
rect 330 440 410 470
rect 470 467 497 513
rect 543 467 600 513
rect 470 440 600 467
rect 180 380 240 440
rect 350 380 410 440
rect 540 380 600 440
rect 180 160 240 210
rect 350 160 410 210
rect 540 160 600 210
<< polycontact >>
rect 357 597 403 643
rect 147 467 193 513
rect 497 467 543 513
<< metal1 >>
rect 0 1198 800 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 800 1198
rect 0 1130 800 1152
rect 130 1007 180 1130
rect 130 773 132 1007
rect 178 773 180 1007
rect 130 720 180 773
rect 420 1000 490 1060
rect 420 860 432 1000
rect 478 860 490 1000
rect 610 1008 660 1130
rect 610 962 612 1008
rect 658 962 660 1008
rect 610 910 660 962
rect 420 780 490 860
rect 420 776 700 780
rect 420 724 624 776
rect 676 724 700 776
rect 420 720 700 724
rect 620 710 690 720
rect 330 646 430 650
rect 330 594 354 646
rect 406 594 430 646
rect 330 590 430 594
rect 120 516 220 520
rect 120 464 144 516
rect 196 464 220 516
rect 120 460 220 464
rect 470 516 570 520
rect 470 464 494 516
rect 546 464 570 516
rect 470 460 570 464
rect 100 350 510 400
rect 100 288 150 350
rect 100 242 102 288
rect 148 242 150 288
rect 100 210 150 242
rect 270 278 320 300
rect 270 232 272 278
rect 318 232 320 278
rect 270 140 320 232
rect 440 288 510 350
rect 440 242 452 288
rect 498 242 510 288
rect 440 210 510 242
rect 630 308 680 710
rect 630 262 632 308
rect 678 262 680 308
rect 630 210 680 262
rect 0 118 800 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 800 118
rect 0 0 800 72
<< via1 >>
rect 624 724 676 776
rect 354 643 406 646
rect 354 597 357 643
rect 357 597 403 643
rect 403 597 406 643
rect 354 594 406 597
rect 144 513 196 516
rect 144 467 147 513
rect 147 467 193 513
rect 193 467 196 513
rect 144 464 196 467
rect 494 513 546 516
rect 494 467 497 513
rect 497 467 543 513
rect 543 467 546 513
rect 494 464 546 467
<< metal2 >>
rect 610 780 690 790
rect 600 776 700 780
rect 600 724 624 776
rect 676 724 700 776
rect 600 720 700 724
rect 610 710 690 720
rect 330 646 430 660
rect 330 594 354 646
rect 406 594 430 646
rect 330 580 430 594
rect 120 516 220 530
rect 120 464 144 516
rect 196 464 220 516
rect 120 450 220 464
rect 470 516 570 530
rect 470 464 494 516
rect 546 464 570 516
rect 470 450 570 464
<< labels >>
rlabel via1 s 144 464 196 516 4 A0
port 1 nsew signal input
rlabel via1 s 354 594 406 646 4 A1
port 2 nsew signal input
rlabel via1 s 494 464 546 516 4 B
port 3 nsew signal input
rlabel via1 s 624 724 676 776 4 Y
port 4 nsew signal output
rlabel metal1 s 130 720 180 1270 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 270 0 320 300 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 610 910 660 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1130 800 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 0 800 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 120 450 220 530 1 A0
port 1 nsew signal input
rlabel metal1 s 120 460 220 520 1 A0
port 1 nsew signal input
rlabel metal2 s 330 580 430 660 1 A1
port 2 nsew signal input
rlabel metal1 s 330 590 430 650 1 A1
port 2 nsew signal input
rlabel metal2 s 470 450 570 530 1 B
port 3 nsew signal input
rlabel metal1 s 470 460 570 520 1 B
port 3 nsew signal input
rlabel metal2 s 610 710 690 790 1 Y
port 4 nsew signal output
rlabel metal2 s 600 720 700 780 1 Y
port 4 nsew signal output
rlabel metal1 s 420 720 490 1060 1 Y
port 4 nsew signal output
rlabel metal1 s 630 210 680 780 1 Y
port 4 nsew signal output
rlabel metal1 s 620 710 690 780 1 Y
port 4 nsew signal output
rlabel metal1 s 420 720 700 780 1 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 800 1270
string GDS_END 342282
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 336862
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
