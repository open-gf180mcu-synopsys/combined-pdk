magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 620 1140 1260
<< nmos >>
rect 200 200 260 370
rect 370 200 430 370
rect 540 200 600 370
rect 710 200 770 370
rect 880 200 940 370
<< pmos >>
rect 200 710 260 1050
rect 370 710 430 1050
rect 540 710 600 1050
rect 710 710 770 1050
rect 880 710 940 1050
<< ndiff >>
rect 100 308 200 370
rect 100 262 122 308
rect 168 262 200 308
rect 100 200 200 262
rect 260 308 370 370
rect 260 262 292 308
rect 338 262 370 308
rect 260 200 370 262
rect 430 308 540 370
rect 430 262 462 308
rect 508 262 540 308
rect 430 200 540 262
rect 600 308 710 370
rect 600 262 632 308
rect 678 262 710 308
rect 600 200 710 262
rect 770 308 880 370
rect 770 262 802 308
rect 848 262 880 308
rect 770 200 880 262
rect 940 308 1040 370
rect 940 262 972 308
rect 1018 262 1040 308
rect 940 200 1040 262
<< pdiff >>
rect 100 997 200 1050
rect 100 763 122 997
rect 168 763 200 997
rect 100 710 200 763
rect 260 997 370 1050
rect 260 763 292 997
rect 338 763 370 997
rect 260 710 370 763
rect 430 1022 540 1050
rect 430 788 462 1022
rect 508 788 540 1022
rect 430 710 540 788
rect 600 997 710 1050
rect 600 763 632 997
rect 678 763 710 997
rect 600 710 710 763
rect 770 1022 880 1050
rect 770 788 802 1022
rect 848 788 880 1022
rect 770 710 880 788
rect 940 997 1040 1050
rect 940 763 972 997
rect 1018 763 1040 997
rect 940 710 1040 763
<< ndiffc >>
rect 122 262 168 308
rect 292 262 338 308
rect 462 262 508 308
rect 632 262 678 308
rect 802 262 848 308
rect 972 262 1018 308
<< pdiffc >>
rect 122 763 168 997
rect 292 763 338 997
rect 462 788 508 1022
rect 632 763 678 997
rect 802 788 848 1022
rect 972 763 1018 997
<< psubdiff >>
rect 70 108 220 130
rect 70 62 122 108
rect 168 62 220 108
rect 70 40 220 62
rect 310 108 460 130
rect 310 62 362 108
rect 408 62 460 108
rect 310 40 460 62
rect 550 108 700 130
rect 550 62 602 108
rect 648 62 700 108
rect 550 40 700 62
rect 790 108 940 130
rect 790 62 842 108
rect 888 62 940 108
rect 790 40 940 62
<< nsubdiff >>
rect 70 1188 220 1210
rect 70 1142 122 1188
rect 168 1142 220 1188
rect 70 1120 220 1142
rect 310 1188 460 1210
rect 310 1142 362 1188
rect 408 1142 460 1188
rect 310 1120 460 1142
rect 550 1188 700 1210
rect 550 1142 602 1188
rect 648 1142 700 1188
rect 550 1120 700 1142
rect 790 1188 940 1210
rect 790 1142 842 1188
rect 888 1142 940 1188
rect 790 1120 940 1142
<< psubdiffcont >>
rect 122 62 168 108
rect 362 62 408 108
rect 602 62 648 108
rect 842 62 888 108
<< nsubdiffcont >>
rect 122 1142 168 1188
rect 362 1142 408 1188
rect 602 1142 648 1188
rect 842 1142 888 1188
<< polysilicon >>
rect 200 1050 260 1100
rect 370 1050 430 1100
rect 540 1050 600 1100
rect 710 1050 770 1100
rect 880 1050 940 1100
rect 200 530 260 710
rect 370 690 430 710
rect 540 690 600 710
rect 710 690 770 710
rect 880 690 940 710
rect 370 680 940 690
rect 310 653 940 680
rect 310 607 337 653
rect 383 630 940 653
rect 383 607 430 630
rect 310 580 430 607
rect 200 503 320 530
rect 200 457 247 503
rect 293 457 320 503
rect 200 430 320 457
rect 370 450 430 580
rect 710 450 770 630
rect 200 370 260 430
rect 370 390 940 450
rect 370 370 430 390
rect 540 370 600 390
rect 710 370 770 390
rect 880 370 940 390
rect 200 150 260 200
rect 370 150 430 200
rect 540 150 600 200
rect 710 150 770 200
rect 880 150 940 200
<< polycontact >>
rect 337 607 383 653
rect 247 457 293 503
<< metal1 >>
rect 0 1188 1140 1260
rect 0 1142 122 1188
rect 168 1142 362 1188
rect 408 1142 602 1188
rect 648 1142 842 1188
rect 888 1142 1140 1188
rect 0 1120 1140 1142
rect 120 997 170 1050
rect 120 763 122 997
rect 168 763 170 997
rect 120 660 170 763
rect 290 997 340 1120
rect 290 763 292 997
rect 338 763 340 997
rect 290 710 340 763
rect 460 1022 510 1050
rect 460 788 462 1022
rect 508 788 510 1022
rect 460 660 510 788
rect 630 997 680 1120
rect 630 763 632 997
rect 678 763 680 997
rect 800 1022 850 1050
rect 800 788 802 1022
rect 848 788 850 1022
rect 800 770 850 788
rect 970 997 1020 1120
rect 630 710 680 763
rect 780 766 880 770
rect 780 714 804 766
rect 856 714 880 766
rect 780 710 880 714
rect 970 763 972 997
rect 1018 763 1020 997
rect 970 710 1020 763
rect 800 660 850 710
rect 120 653 410 660
rect 120 607 337 653
rect 383 607 410 653
rect 120 600 410 607
rect 460 600 850 660
rect 120 308 170 600
rect 220 506 320 510
rect 220 454 244 506
rect 296 454 320 506
rect 220 450 320 454
rect 460 480 510 600
rect 800 480 850 600
rect 460 420 850 480
rect 120 262 122 308
rect 168 262 170 308
rect 120 200 170 262
rect 290 308 340 370
rect 290 262 292 308
rect 338 262 340 308
rect 290 130 340 262
rect 460 308 510 420
rect 460 262 462 308
rect 508 262 510 308
rect 460 200 510 262
rect 630 308 680 370
rect 630 262 632 308
rect 678 262 680 308
rect 630 130 680 262
rect 800 308 850 420
rect 800 262 802 308
rect 848 262 850 308
rect 800 200 850 262
rect 970 308 1020 370
rect 970 262 972 308
rect 1018 262 1020 308
rect 970 130 1020 262
rect 0 108 1140 130
rect 0 62 122 108
rect 168 62 362 108
rect 408 62 602 108
rect 648 62 842 108
rect 888 62 1140 108
rect 0 -10 1140 62
<< via1 >>
rect 804 714 856 766
rect 244 503 296 506
rect 244 457 247 503
rect 247 457 293 503
rect 293 457 296 503
rect 244 454 296 457
<< metal2 >>
rect 780 766 880 780
rect 780 714 804 766
rect 856 714 880 766
rect 780 700 880 714
rect 230 510 310 520
rect 220 506 320 510
rect 220 454 244 506
rect 296 454 320 506
rect 220 450 320 454
rect 230 440 310 450
<< labels >>
rlabel via1 s 244 454 296 506 4 A
port 1 nsew signal input
rlabel via1 s 804 714 856 766 4 Y
port 2 nsew signal output
rlabel metal1 s 290 710 340 1260 4 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 290 -10 340 370 4 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 630 710 680 1260 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 970 710 1020 1260 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 1120 1140 1260 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 630 -10 680 370 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 970 -10 1020 370 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -10 1140 130 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal2 s 230 440 310 520 1 A
port 1 nsew signal input
rlabel metal2 s 220 450 320 510 1 A
port 1 nsew signal input
rlabel metal1 s 220 450 320 510 1 A
port 1 nsew signal input
rlabel metal2 s 780 700 880 780 1 Y
port 2 nsew signal output
rlabel metal1 s 460 200 510 1050 1 Y
port 2 nsew signal output
rlabel metal1 s 460 420 850 480 1 Y
port 2 nsew signal output
rlabel metal1 s 460 600 850 660 1 Y
port 2 nsew signal output
rlabel metal1 s 800 200 850 1050 1 Y
port 2 nsew signal output
rlabel metal1 s 780 710 880 770 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -10 1140 1260
string GDS_END 111746
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 104930
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
