magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 565 390 635
rect 140 435 165 565
rect 310 390 335 530
rect 300 388 350 390
rect 300 362 312 388
rect 338 362 350 388
rect 300 360 350 362
rect 160 323 210 325
rect 160 297 172 323
rect 198 297 210 323
rect 160 295 210 297
rect 60 258 110 260
rect 60 232 72 258
rect 98 232 110 258
rect 60 230 110 232
rect 235 258 285 260
rect 235 232 247 258
rect 273 232 285 258
rect 235 230 285 232
rect 310 200 335 360
rect 70 70 95 190
rect 210 175 335 200
rect 210 105 235 175
rect 295 70 320 150
rect 0 0 390 70
<< via1 >>
rect 312 362 338 388
rect 172 297 198 323
rect 72 232 98 258
rect 247 232 273 258
<< obsm1 >>
rect 55 410 80 530
rect 225 410 250 530
rect 55 385 250 410
<< metal2 >>
rect 300 388 350 395
rect 300 362 312 388
rect 338 362 350 388
rect 300 355 350 362
rect 160 323 210 330
rect 160 297 172 323
rect 198 297 210 323
rect 160 290 210 297
rect 60 258 110 265
rect 60 232 72 258
rect 98 232 110 258
rect 60 225 110 232
rect 235 258 285 265
rect 235 232 247 258
rect 273 232 285 258
rect 235 225 285 232
<< labels >>
rlabel metal1 s 140 435 165 635 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 565 390 635 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 70 0 95 190 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 295 0 320 150 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 390 70 6 VSS
port 6 nsew ground bidirectional abutment
rlabel via1 s 72 232 98 258 6 A0
port 2 nsew signal input
rlabel metal2 s 60 225 110 265 6 A0
port 2 nsew signal input
rlabel metal1 s 60 230 110 260 6 A0
port 2 nsew signal input
rlabel via1 s 172 297 198 323 6 A1
port 3 nsew signal input
rlabel metal2 s 160 290 210 330 6 A1
port 3 nsew signal input
rlabel metal1 s 160 295 210 325 6 A1
port 3 nsew signal input
rlabel via1 s 247 232 273 258 6 B
port 4 nsew signal input
rlabel metal2 s 235 225 285 265 6 B
port 4 nsew signal input
rlabel metal1 s 235 230 285 260 6 B
port 4 nsew signal input
rlabel via1 s 312 362 338 388 6 Y
port 1 nsew signal output
rlabel metal2 s 300 355 350 395 6 Y
port 1 nsew signal output
rlabel metal1 s 210 105 235 200 6 Y
port 1 nsew signal output
rlabel metal1 s 210 175 335 200 6 Y
port 1 nsew signal output
rlabel metal1 s 310 175 335 530 6 Y
port 1 nsew signal output
rlabel metal1 s 300 360 350 390 6 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 390 635
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 46002
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 40774
<< end >>
