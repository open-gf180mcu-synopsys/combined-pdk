magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 1878 870
<< pwell >>
rect -86 -86 1878 352
<< metal1 >>
rect 0 724 1792 844
rect 297 657 365 724
rect 1313 635 1381 724
rect 1643 542 1720 639
rect 1362 466 1720 542
rect 186 240 671 320
rect 317 60 385 127
rect 1344 60 1390 138
rect 1674 135 1720 466
rect 0 -60 1792 60
<< obsm1 >>
rect 49 481 117 621
rect 49 413 653 481
rect 49 180 95 413
rect 744 382 790 632
rect 908 493 954 632
rect 908 447 1231 493
rect 744 336 1097 382
rect 49 134 117 180
rect 744 154 821 336
rect 1167 325 1231 447
rect 1167 279 1595 325
rect 1167 211 1231 279
rect 908 143 1231 211
<< labels >>
rlabel metal1 s 186 240 671 320 6 I
port 1 nsew default input
rlabel metal1 s 1674 135 1720 466 6 Z
port 2 nsew default output
rlabel metal1 s 1362 466 1720 542 6 Z
port 2 nsew default output
rlabel metal1 s 1643 542 1720 639 6 Z
port 2 nsew default output
rlabel metal1 s 1313 635 1381 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 1792 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 1878 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 1878 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 1792 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1344 60 1390 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1094044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1090088
<< end >>
