magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 780 1660
<< nmos >>
rect 180 210 240 380
rect 350 210 410 380
rect 520 210 580 380
<< pmos >>
rect 210 1110 270 1450
rect 330 1110 390 1450
rect 500 1110 560 1450
<< ndiff >>
rect 80 318 180 380
rect 80 272 102 318
rect 148 272 180 318
rect 80 210 180 272
rect 240 288 350 380
rect 240 242 272 288
rect 318 242 350 288
rect 240 210 350 242
rect 410 318 520 380
rect 410 272 442 318
rect 488 272 520 318
rect 410 210 520 272
rect 580 318 680 380
rect 580 272 612 318
rect 658 272 680 318
rect 580 210 680 272
<< pdiff >>
rect 110 1397 210 1450
rect 110 1163 132 1397
rect 178 1163 210 1397
rect 110 1110 210 1163
rect 270 1110 330 1450
rect 390 1397 500 1450
rect 390 1163 422 1397
rect 468 1163 500 1397
rect 390 1110 500 1163
rect 560 1397 660 1450
rect 560 1163 592 1397
rect 638 1163 660 1397
rect 560 1110 660 1163
<< ndiffc >>
rect 102 272 148 318
rect 272 242 318 288
rect 442 272 488 318
rect 612 272 658 318
<< pdiffc >>
rect 132 1163 178 1397
rect 422 1163 468 1397
rect 592 1163 638 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
<< polysilicon >>
rect 210 1450 270 1500
rect 330 1450 390 1500
rect 500 1450 560 1500
rect 210 1090 270 1110
rect 160 1050 270 1090
rect 160 800 220 1050
rect 330 930 390 1110
rect 270 903 390 930
rect 270 857 317 903
rect 363 857 390 903
rect 270 830 390 857
rect 80 773 220 800
rect 80 727 117 773
rect 163 727 220 773
rect 80 700 220 727
rect 160 470 220 700
rect 330 470 390 830
rect 500 800 560 1110
rect 440 773 560 800
rect 440 727 467 773
rect 513 727 560 773
rect 440 700 560 727
rect 500 470 560 700
rect 160 440 240 470
rect 330 440 410 470
rect 500 440 580 470
rect 180 380 240 440
rect 350 380 410 440
rect 520 380 580 440
rect 180 160 240 210
rect 350 160 410 210
rect 520 160 580 210
<< polycontact >>
rect 317 857 363 903
rect 117 727 163 773
rect 467 727 513 773
<< metal1 >>
rect 0 1588 780 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 780 1588
rect 0 1520 780 1542
rect 130 1397 180 1520
rect 130 1163 132 1397
rect 178 1163 180 1397
rect 130 1110 180 1163
rect 420 1397 470 1450
rect 420 1163 422 1397
rect 468 1163 470 1397
rect 420 1040 470 1163
rect 590 1397 640 1520
rect 590 1163 592 1397
rect 638 1163 640 1397
rect 590 1110 640 1163
rect 420 1036 670 1040
rect 420 984 594 1036
rect 646 984 670 1036
rect 420 980 670 984
rect 290 906 390 910
rect 290 854 314 906
rect 366 854 390 906
rect 290 850 390 854
rect 90 776 190 780
rect 90 724 114 776
rect 166 724 190 776
rect 90 720 190 724
rect 440 776 540 780
rect 440 724 464 776
rect 516 724 540 776
rect 440 720 540 724
rect 590 520 640 980
rect 590 470 660 520
rect 100 370 490 420
rect 100 318 150 370
rect 100 272 102 318
rect 148 272 150 318
rect 100 210 150 272
rect 270 288 320 320
rect 270 242 272 288
rect 318 242 320 288
rect 270 140 320 242
rect 440 318 490 370
rect 440 272 442 318
rect 488 272 490 318
rect 440 210 490 272
rect 610 318 660 470
rect 610 272 612 318
rect 658 272 660 318
rect 610 210 660 272
rect 0 118 780 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 780 118
rect 0 0 780 72
<< via1 >>
rect 594 984 646 1036
rect 314 903 366 906
rect 314 857 317 903
rect 317 857 363 903
rect 363 857 366 903
rect 314 854 366 857
rect 114 773 166 776
rect 114 727 117 773
rect 117 727 163 773
rect 163 727 166 773
rect 114 724 166 727
rect 464 773 516 776
rect 464 727 467 773
rect 467 727 513 773
rect 513 727 516 773
rect 464 724 516 727
<< metal2 >>
rect 570 1036 670 1050
rect 570 984 594 1036
rect 646 984 670 1036
rect 570 970 670 984
rect 290 906 390 920
rect 290 854 314 906
rect 366 854 390 906
rect 290 840 390 854
rect 90 776 190 790
rect 90 724 114 776
rect 166 724 190 776
rect 90 710 190 724
rect 440 776 540 790
rect 440 724 464 776
rect 516 724 540 776
rect 440 710 540 724
<< labels >>
rlabel via1 s 114 724 166 776 4 A0
port 1 nsew signal input
rlabel via1 s 314 854 366 906 4 A1
port 2 nsew signal input
rlabel via1 s 464 724 516 776 4 B
port 3 nsew signal input
rlabel via1 s 594 984 646 1036 4 Y
port 4 nsew signal output
rlabel metal1 s 130 1110 180 1660 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 270 0 320 320 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 590 1110 640 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1520 780 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 0 780 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 90 710 190 790 1 A0
port 1 nsew signal input
rlabel metal1 s 90 720 190 780 1 A0
port 1 nsew signal input
rlabel metal2 s 290 840 390 920 1 A1
port 2 nsew signal input
rlabel metal1 s 290 850 390 910 1 A1
port 2 nsew signal input
rlabel metal2 s 440 710 540 790 1 B
port 3 nsew signal input
rlabel metal1 s 440 720 540 780 1 B
port 3 nsew signal input
rlabel metal2 s 570 970 670 1050 1 Y
port 4 nsew signal output
rlabel metal1 s 420 980 470 1450 1 Y
port 4 nsew signal output
rlabel metal1 s 590 470 640 1040 1 Y
port 4 nsew signal output
rlabel metal1 s 610 210 660 520 1 Y
port 4 nsew signal output
rlabel metal1 s 420 980 670 1040 1 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 780 1660
string GDS_END 478352
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 472740
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
