magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3850 1660
<< nmos >>
rect 190 210 250 380
rect 540 210 600 380
rect 710 210 770 380
rect 1060 210 1120 380
rect 1220 210 1280 380
rect 1390 210 1450 380
rect 1500 210 1560 380
rect 1670 210 1730 380
rect 1780 210 1840 380
rect 1950 210 2010 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2590 210 2650 380
rect 2910 210 2970 380
rect 3080 210 3140 380
rect 3430 210 3490 380
rect 3600 210 3660 380
<< pmos >>
rect 190 1110 250 1450
rect 510 1110 570 1450
rect 620 1110 680 1450
rect 1060 1110 1120 1450
rect 1220 1110 1280 1450
rect 1390 1110 1450 1450
rect 1500 1110 1560 1450
rect 1670 1110 1730 1450
rect 1780 1110 1840 1450
rect 1950 1110 2010 1450
rect 2060 1110 2120 1450
rect 2230 1110 2290 1450
rect 2590 1110 2650 1450
rect 3000 1110 3060 1450
rect 3110 1110 3170 1450
rect 3430 1110 3490 1450
rect 3600 1110 3660 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 440 318 540 380
rect 440 272 462 318
rect 508 272 540 318
rect 440 210 540 272
rect 600 318 710 380
rect 600 272 632 318
rect 678 272 710 318
rect 600 210 710 272
rect 770 318 870 380
rect 770 272 802 318
rect 848 272 870 318
rect 770 210 870 272
rect 960 318 1060 380
rect 960 272 982 318
rect 1028 272 1060 318
rect 960 210 1060 272
rect 1120 210 1220 380
rect 1280 318 1390 380
rect 1280 272 1312 318
rect 1358 272 1390 318
rect 1280 210 1390 272
rect 1450 210 1500 380
rect 1560 278 1670 380
rect 1560 232 1592 278
rect 1638 232 1670 278
rect 1560 210 1670 232
rect 1730 210 1780 380
rect 1840 318 1950 380
rect 1840 272 1872 318
rect 1918 272 1950 318
rect 1840 210 1950 272
rect 2010 210 2060 380
rect 2120 318 2230 380
rect 2120 272 2152 318
rect 2198 272 2230 318
rect 2120 210 2230 272
rect 2290 318 2390 380
rect 2290 272 2322 318
rect 2368 272 2390 318
rect 2290 210 2390 272
rect 2490 318 2590 380
rect 2490 272 2512 318
rect 2558 272 2590 318
rect 2490 210 2590 272
rect 2650 318 2750 380
rect 2650 272 2682 318
rect 2728 272 2750 318
rect 2650 210 2750 272
rect 2810 318 2910 380
rect 2810 272 2832 318
rect 2878 272 2910 318
rect 2810 210 2910 272
rect 2970 318 3080 380
rect 2970 272 3002 318
rect 3048 272 3080 318
rect 2970 210 3080 272
rect 3140 318 3240 380
rect 3140 272 3172 318
rect 3218 272 3240 318
rect 3140 210 3240 272
rect 3330 318 3430 380
rect 3330 272 3352 318
rect 3398 272 3430 318
rect 3330 210 3430 272
rect 3490 318 3600 380
rect 3490 272 3522 318
rect 3568 272 3600 318
rect 3490 210 3600 272
rect 3660 318 3760 380
rect 3660 272 3692 318
rect 3738 272 3760 318
rect 3660 210 3760 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 350 1450
rect 250 1163 282 1397
rect 328 1163 350 1397
rect 250 1110 350 1163
rect 410 1397 510 1450
rect 410 1163 432 1397
rect 478 1163 510 1397
rect 410 1110 510 1163
rect 570 1110 620 1450
rect 680 1397 780 1450
rect 680 1163 712 1397
rect 758 1163 780 1397
rect 680 1110 780 1163
rect 960 1397 1060 1450
rect 960 1163 982 1397
rect 1028 1163 1060 1397
rect 960 1110 1060 1163
rect 1120 1110 1220 1450
rect 1280 1397 1390 1450
rect 1280 1163 1312 1397
rect 1358 1163 1390 1397
rect 1280 1110 1390 1163
rect 1450 1110 1500 1450
rect 1560 1397 1670 1450
rect 1560 1163 1592 1397
rect 1638 1163 1670 1397
rect 1560 1110 1670 1163
rect 1730 1110 1780 1450
rect 1840 1425 1950 1450
rect 1840 1285 1872 1425
rect 1918 1285 1950 1425
rect 1840 1110 1950 1285
rect 2010 1110 2060 1450
rect 2120 1425 2230 1450
rect 2120 1285 2152 1425
rect 2198 1285 2230 1425
rect 2120 1110 2230 1285
rect 2290 1397 2390 1450
rect 2290 1163 2322 1397
rect 2368 1163 2390 1397
rect 2290 1110 2390 1163
rect 2490 1397 2590 1450
rect 2490 1163 2512 1397
rect 2558 1163 2590 1397
rect 2490 1110 2590 1163
rect 2650 1397 2750 1450
rect 2650 1163 2682 1397
rect 2728 1163 2750 1397
rect 2650 1110 2750 1163
rect 2900 1397 3000 1450
rect 2900 1163 2922 1397
rect 2968 1163 3000 1397
rect 2900 1110 3000 1163
rect 3060 1110 3110 1450
rect 3170 1397 3270 1450
rect 3170 1163 3202 1397
rect 3248 1163 3270 1397
rect 3170 1110 3270 1163
rect 3330 1397 3430 1450
rect 3330 1163 3352 1397
rect 3398 1163 3430 1397
rect 3330 1110 3430 1163
rect 3490 1397 3600 1450
rect 3490 1163 3522 1397
rect 3568 1163 3600 1397
rect 3490 1110 3600 1163
rect 3660 1397 3760 1450
rect 3660 1163 3692 1397
rect 3738 1163 3760 1397
rect 3660 1110 3760 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 462 272 508 318
rect 632 272 678 318
rect 802 272 848 318
rect 982 272 1028 318
rect 1312 272 1358 318
rect 1592 232 1638 278
rect 1872 272 1918 318
rect 2152 272 2198 318
rect 2322 272 2368 318
rect 2512 272 2558 318
rect 2682 272 2728 318
rect 2832 272 2878 318
rect 3002 272 3048 318
rect 3172 272 3218 318
rect 3352 272 3398 318
rect 3522 272 3568 318
rect 3692 272 3738 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 432 1163 478 1397
rect 712 1163 758 1397
rect 982 1163 1028 1397
rect 1312 1163 1358 1397
rect 1592 1163 1638 1397
rect 1872 1285 1918 1425
rect 2152 1285 2198 1425
rect 2322 1163 2368 1397
rect 2512 1163 2558 1397
rect 2682 1163 2728 1397
rect 2922 1163 2968 1397
rect 3202 1163 3248 1397
rect 3352 1163 3398 1397
rect 3522 1163 3568 1397
rect 3692 1163 3738 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
rect 980 118 1130 140
rect 980 72 1032 118
rect 1078 72 1130 118
rect 980 50 1130 72
rect 1210 118 1360 140
rect 1210 72 1262 118
rect 1308 72 1360 118
rect 1210 50 1360 72
rect 1440 118 1590 140
rect 1440 72 1492 118
rect 1538 72 1590 118
rect 1440 50 1590 72
rect 1670 118 1820 140
rect 1670 72 1722 118
rect 1768 72 1820 118
rect 1670 50 1820 72
rect 1900 118 2050 140
rect 1900 72 1952 118
rect 1998 72 2050 118
rect 1900 50 2050 72
rect 2130 118 2280 140
rect 2130 72 2182 118
rect 2228 72 2280 118
rect 2130 50 2280 72
rect 2360 118 2510 140
rect 2360 72 2412 118
rect 2458 72 2510 118
rect 2360 50 2510 72
rect 2590 118 2740 140
rect 2590 72 2642 118
rect 2688 72 2740 118
rect 2590 50 2740 72
rect 2820 118 2970 140
rect 2820 72 2872 118
rect 2918 72 2970 118
rect 2820 50 2970 72
rect 3050 118 3200 140
rect 3050 72 3102 118
rect 3148 72 3200 118
rect 3050 50 3200 72
rect 3280 118 3430 140
rect 3280 72 3332 118
rect 3378 72 3430 118
rect 3280 50 3430 72
rect 3510 118 3660 140
rect 3510 72 3562 118
rect 3608 72 3660 118
rect 3510 50 3660 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
rect 980 1588 1130 1610
rect 980 1542 1032 1588
rect 1078 1542 1130 1588
rect 980 1520 1130 1542
rect 1210 1588 1360 1610
rect 1210 1542 1262 1588
rect 1308 1542 1360 1588
rect 1210 1520 1360 1542
rect 1440 1588 1590 1610
rect 1440 1542 1492 1588
rect 1538 1542 1590 1588
rect 1440 1520 1590 1542
rect 1670 1588 1820 1610
rect 1670 1542 1722 1588
rect 1768 1542 1820 1588
rect 1670 1520 1820 1542
rect 1900 1588 2050 1610
rect 1900 1542 1952 1588
rect 1998 1542 2050 1588
rect 1900 1520 2050 1542
rect 2130 1588 2280 1610
rect 2130 1542 2182 1588
rect 2228 1542 2280 1588
rect 2130 1520 2280 1542
rect 2360 1588 2510 1610
rect 2360 1542 2412 1588
rect 2458 1542 2510 1588
rect 2360 1520 2510 1542
rect 2590 1588 2740 1610
rect 2590 1542 2642 1588
rect 2688 1542 2740 1588
rect 2590 1520 2740 1542
rect 2820 1588 2970 1610
rect 2820 1542 2872 1588
rect 2918 1542 2970 1588
rect 2820 1520 2970 1542
rect 3050 1588 3200 1610
rect 3050 1542 3102 1588
rect 3148 1542 3200 1588
rect 3050 1520 3200 1542
rect 3280 1588 3430 1610
rect 3280 1542 3332 1588
rect 3378 1542 3430 1588
rect 3280 1520 3430 1542
rect 3510 1588 3660 1610
rect 3510 1542 3562 1588
rect 3608 1542 3660 1588
rect 3510 1520 3660 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
rect 1032 72 1078 118
rect 1262 72 1308 118
rect 1492 72 1538 118
rect 1722 72 1768 118
rect 1952 72 1998 118
rect 2182 72 2228 118
rect 2412 72 2458 118
rect 2642 72 2688 118
rect 2872 72 2918 118
rect 3102 72 3148 118
rect 3332 72 3378 118
rect 3562 72 3608 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
rect 1032 1542 1078 1588
rect 1262 1542 1308 1588
rect 1492 1542 1538 1588
rect 1722 1542 1768 1588
rect 1952 1542 1998 1588
rect 2182 1542 2228 1588
rect 2412 1542 2458 1588
rect 2642 1542 2688 1588
rect 2872 1542 2918 1588
rect 3102 1542 3148 1588
rect 3332 1542 3378 1588
rect 3562 1542 3608 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 510 1450 570 1500
rect 620 1450 680 1500
rect 1060 1450 1120 1500
rect 1220 1450 1280 1500
rect 1390 1450 1450 1500
rect 1500 1450 1560 1500
rect 1670 1450 1730 1500
rect 1780 1450 1840 1500
rect 1950 1450 2010 1500
rect 2060 1450 2120 1500
rect 2230 1450 2290 1500
rect 2590 1450 2650 1500
rect 3000 1450 3060 1500
rect 3110 1450 3170 1500
rect 3430 1450 3490 1500
rect 3600 1450 3660 1500
rect 190 1060 250 1110
rect 120 1038 250 1060
rect 120 992 142 1038
rect 188 992 250 1038
rect 120 970 250 992
rect 190 380 250 970
rect 510 800 570 1110
rect 620 1060 680 1110
rect 620 1000 770 1060
rect 710 930 770 1000
rect 710 903 880 930
rect 710 857 797 903
rect 843 857 880 903
rect 710 830 880 857
rect 510 773 630 800
rect 510 727 557 773
rect 603 727 630 773
rect 510 700 630 727
rect 510 650 570 700
rect 510 610 600 650
rect 540 380 600 610
rect 710 380 770 830
rect 1060 800 1120 1110
rect 1220 930 1280 1110
rect 1220 903 1320 930
rect 1220 857 1247 903
rect 1293 857 1320 903
rect 1220 830 1320 857
rect 1060 773 1180 800
rect 1060 727 1107 773
rect 1153 727 1180 773
rect 1060 700 1180 727
rect 1060 380 1120 700
rect 1390 660 1450 1110
rect 1500 1060 1560 1110
rect 1670 1060 1730 1110
rect 1500 1033 1730 1060
rect 1500 990 1537 1033
rect 1510 987 1537 990
rect 1583 990 1730 1033
rect 1583 987 1610 990
rect 1510 940 1610 987
rect 1780 660 1840 1110
rect 1950 930 2010 1110
rect 1910 903 2010 930
rect 1910 857 1937 903
rect 1983 857 2010 903
rect 1910 830 2010 857
rect 2060 800 2120 1110
rect 2230 930 2290 1110
rect 2230 903 2330 930
rect 2230 857 2257 903
rect 2303 857 2330 903
rect 2230 830 2330 857
rect 2050 773 2150 800
rect 2050 727 2077 773
rect 2123 727 2150 773
rect 2050 700 2150 727
rect 1910 660 2010 670
rect 1220 643 2010 660
rect 1220 600 1937 643
rect 1220 380 1280 600
rect 1910 597 1937 600
rect 1983 597 2010 643
rect 1910 570 2010 597
rect 1350 513 1450 540
rect 1510 520 1610 540
rect 1350 467 1377 513
rect 1423 467 1450 513
rect 1350 440 1450 467
rect 1390 380 1450 440
rect 1500 513 1730 520
rect 1500 467 1537 513
rect 1583 467 1730 513
rect 1500 440 1730 467
rect 1500 380 1560 440
rect 1670 380 1730 440
rect 1780 503 1880 530
rect 1780 457 1807 503
rect 1853 457 1880 503
rect 1780 430 1880 457
rect 1780 380 1840 430
rect 1950 380 2010 570
rect 2060 380 2120 700
rect 2230 380 2290 830
rect 2590 670 2650 1110
rect 3000 1060 3060 1110
rect 2880 1000 3060 1060
rect 2590 648 2720 670
rect 2590 602 2652 648
rect 2698 602 2720 648
rect 2590 580 2720 602
rect 2590 380 2650 580
rect 2880 530 2940 1000
rect 3110 650 3170 1110
rect 3430 670 3490 1110
rect 3600 930 3660 1110
rect 3540 903 3660 930
rect 3540 857 3567 903
rect 3613 857 3660 903
rect 3540 830 3660 857
rect 2800 503 2940 530
rect 2800 457 2837 503
rect 2883 470 2940 503
rect 3080 610 3170 650
rect 3370 643 3490 670
rect 3080 530 3140 610
rect 3370 597 3417 643
rect 3463 597 3490 643
rect 3370 570 3490 597
rect 3080 503 3200 530
rect 2883 457 2970 470
rect 2800 430 2970 457
rect 2910 380 2970 430
rect 3080 457 3127 503
rect 3173 457 3200 503
rect 3080 430 3200 457
rect 3080 380 3140 430
rect 3430 380 3490 570
rect 3600 380 3660 830
rect 190 160 250 210
rect 540 160 600 210
rect 710 160 770 210
rect 1060 160 1120 210
rect 1220 160 1280 210
rect 1390 160 1450 210
rect 1500 160 1560 210
rect 1670 160 1730 210
rect 1780 160 1840 210
rect 1950 160 2010 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2590 160 2650 210
rect 2910 160 2970 210
rect 3080 160 3140 210
rect 3430 160 3490 210
rect 3600 160 3660 210
<< polycontact >>
rect 142 992 188 1038
rect 797 857 843 903
rect 557 727 603 773
rect 1247 857 1293 903
rect 1107 727 1153 773
rect 1537 987 1583 1033
rect 1937 857 1983 903
rect 2257 857 2303 903
rect 2077 727 2123 773
rect 1937 597 1983 643
rect 1377 467 1423 513
rect 1537 467 1583 513
rect 1807 457 1853 503
rect 2652 602 2698 648
rect 3567 857 3613 903
rect 2837 457 2883 503
rect 3417 597 3463 643
rect 3127 457 3173 503
<< metal1 >>
rect 0 1588 3850 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1032 1588
rect 1078 1542 1262 1588
rect 1308 1542 1492 1588
rect 1538 1542 1722 1588
rect 1768 1542 1952 1588
rect 1998 1542 2182 1588
rect 2228 1542 2412 1588
rect 2458 1542 2642 1588
rect 2688 1542 2872 1588
rect 2918 1542 3102 1588
rect 3148 1542 3332 1588
rect 3378 1542 3562 1588
rect 3608 1542 3850 1588
rect 0 1520 3850 1542
rect 110 1397 160 1520
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1110 160 1163
rect 280 1397 330 1450
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 110 1038 210 1040
rect 110 1036 142 1038
rect 110 984 134 1036
rect 188 992 210 1038
rect 186 984 210 992
rect 110 980 210 984
rect 280 520 330 1163
rect 430 1397 480 1450
rect 430 1163 432 1397
rect 478 1163 480 1397
rect 430 570 480 1163
rect 710 1397 760 1520
rect 710 1163 712 1397
rect 758 1163 760 1397
rect 710 1110 760 1163
rect 980 1397 1030 1520
rect 980 1163 982 1397
rect 1028 1163 1030 1397
rect 980 1110 1030 1163
rect 1310 1397 1360 1450
rect 1310 1163 1312 1397
rect 1358 1163 1360 1397
rect 1310 1060 1360 1163
rect 1590 1397 1640 1520
rect 1590 1163 1592 1397
rect 1638 1163 1640 1397
rect 1870 1425 1920 1450
rect 1870 1285 1872 1425
rect 1918 1285 1920 1425
rect 1870 1260 1920 1285
rect 2150 1425 2200 1520
rect 2150 1285 2152 1425
rect 2198 1285 2200 1425
rect 2150 1260 2200 1285
rect 2320 1397 2370 1450
rect 1590 1110 1640 1163
rect 1690 1210 1920 1260
rect 980 1010 1360 1060
rect 1510 1033 1610 1040
rect 980 910 1030 1010
rect 1510 987 1537 1033
rect 1583 987 1610 1033
rect 1510 980 1610 987
rect 770 903 1030 910
rect 770 857 797 903
rect 843 857 1030 903
rect 770 850 1030 857
rect 1220 906 1450 910
rect 1220 903 1374 906
rect 1220 857 1247 903
rect 1293 857 1374 903
rect 1220 854 1374 857
rect 1426 854 1450 906
rect 1220 850 1450 854
rect 530 776 630 780
rect 530 724 554 776
rect 606 724 630 776
rect 530 720 630 724
rect 430 520 680 570
rect 790 520 840 530
rect 980 520 1030 850
rect 1080 776 1180 780
rect 1080 724 1104 776
rect 1156 724 1180 776
rect 1080 720 1180 724
rect 1370 520 1430 850
rect 1530 520 1590 980
rect 1690 760 1740 1210
rect 2320 1163 2322 1397
rect 2368 1163 2370 1397
rect 2040 1036 2140 1040
rect 2040 984 2064 1036
rect 2116 984 2140 1036
rect 2040 980 2140 984
rect 2320 1020 2370 1163
rect 2510 1397 2560 1450
rect 2510 1163 2512 1397
rect 2558 1163 2560 1397
rect 1680 710 1740 760
rect 1800 906 2010 910
rect 1800 854 1934 906
rect 1986 854 2010 906
rect 1800 850 2010 854
rect 260 516 360 520
rect 260 464 284 516
rect 336 464 360 516
rect 260 460 360 464
rect 600 516 870 520
rect 600 464 794 516
rect 846 464 870 516
rect 980 470 1180 520
rect 600 460 870 464
rect 280 450 340 460
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 450
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 460 318 510 380
rect 460 272 462 318
rect 508 272 510 318
rect 460 140 510 272
rect 630 318 680 460
rect 790 450 840 460
rect 1100 380 1180 470
rect 1350 513 1450 520
rect 1350 467 1377 513
rect 1423 467 1450 513
rect 1350 460 1450 467
rect 1510 516 1610 520
rect 1510 464 1534 516
rect 1586 464 1610 516
rect 1510 460 1610 464
rect 1680 390 1730 710
rect 1800 510 1860 850
rect 2060 780 2120 980
rect 2320 970 2430 1020
rect 2230 906 2330 910
rect 2230 854 2254 906
rect 2306 854 2330 906
rect 2230 850 2330 854
rect 2380 780 2430 970
rect 2510 910 2560 1163
rect 2680 1397 2730 1520
rect 2680 1163 2682 1397
rect 2728 1163 2730 1397
rect 2680 1110 2730 1163
rect 2920 1397 2970 1520
rect 2920 1163 2922 1397
rect 2968 1163 2970 1397
rect 2920 1110 2970 1163
rect 3200 1397 3250 1450
rect 3200 1163 3202 1397
rect 3248 1163 3250 1397
rect 2830 1040 2890 1060
rect 3200 1040 3250 1163
rect 3350 1397 3400 1450
rect 3350 1163 3352 1397
rect 3398 1163 3400 1397
rect 2830 1036 3280 1040
rect 2830 984 2834 1036
rect 2886 984 3204 1036
rect 3256 984 3280 1036
rect 2830 980 3280 984
rect 2830 960 2890 980
rect 2480 906 2580 910
rect 2480 854 2504 906
rect 2556 854 2580 906
rect 2480 850 2580 854
rect 2050 776 2150 780
rect 2050 724 2074 776
rect 2126 724 2150 776
rect 2050 720 2150 724
rect 2320 730 2430 780
rect 1910 646 2010 650
rect 1910 594 1934 646
rect 1986 594 2010 646
rect 1910 590 2010 594
rect 2320 646 2380 730
rect 2320 594 2324 646
rect 2376 594 2380 646
rect 2320 570 2380 594
rect 1780 503 1880 510
rect 1780 457 1807 503
rect 1853 457 1880 503
rect 1780 450 1880 457
rect 1680 386 1950 390
rect 630 272 632 318
rect 678 272 680 318
rect 630 210 680 272
rect 800 318 850 380
rect 800 272 802 318
rect 848 272 850 318
rect 800 140 850 272
rect 980 318 1030 380
rect 1100 330 1360 380
rect 1680 340 1874 386
rect 980 272 982 318
rect 1028 272 1030 318
rect 980 140 1030 272
rect 1310 318 1360 330
rect 1310 272 1312 318
rect 1358 272 1360 318
rect 1870 334 1874 340
rect 1926 334 1950 386
rect 1870 330 1950 334
rect 1870 318 1920 330
rect 1310 210 1360 272
rect 1590 278 1640 300
rect 1590 232 1592 278
rect 1638 232 1640 278
rect 1590 140 1640 232
rect 1870 272 1872 318
rect 1918 272 1920 318
rect 1870 210 1920 272
rect 2150 318 2200 380
rect 2150 272 2152 318
rect 2198 272 2200 318
rect 2150 140 2200 272
rect 2320 318 2370 570
rect 2320 272 2322 318
rect 2368 272 2370 318
rect 2320 210 2370 272
rect 2510 318 2560 850
rect 3200 650 3250 980
rect 3350 910 3400 1163
rect 3520 1397 3570 1520
rect 3520 1163 3522 1397
rect 3568 1163 3570 1397
rect 3520 1110 3570 1163
rect 3690 1397 3740 1450
rect 3690 1163 3692 1397
rect 3738 1163 3740 1397
rect 3690 1050 3740 1163
rect 3690 1036 3790 1050
rect 3690 984 3714 1036
rect 3766 984 3790 1036
rect 3690 980 3790 984
rect 3690 970 3780 980
rect 3350 906 3640 910
rect 3350 854 3564 906
rect 3616 854 3640 906
rect 3350 850 3640 854
rect 2630 648 2730 650
rect 2630 602 2652 648
rect 2698 646 2730 648
rect 2630 594 2654 602
rect 2706 594 2730 646
rect 2630 590 2730 594
rect 3000 646 3490 650
rect 3000 594 3414 646
rect 3466 594 3490 646
rect 3000 590 3490 594
rect 2810 506 2910 510
rect 2810 454 2834 506
rect 2886 454 2910 506
rect 2810 450 2910 454
rect 2510 272 2512 318
rect 2558 272 2560 318
rect 2510 210 2560 272
rect 2680 318 2730 380
rect 2680 272 2682 318
rect 2728 272 2730 318
rect 2680 140 2730 272
rect 2830 318 2880 380
rect 2830 272 2832 318
rect 2878 272 2880 318
rect 2830 140 2880 272
rect 3000 318 3050 590
rect 3100 506 3200 510
rect 3100 454 3124 506
rect 3176 454 3200 506
rect 3570 480 3620 850
rect 3100 450 3200 454
rect 3350 430 3620 480
rect 3000 272 3002 318
rect 3048 272 3050 318
rect 3000 210 3050 272
rect 3170 318 3220 380
rect 3170 272 3172 318
rect 3218 272 3220 318
rect 3170 140 3220 272
rect 3350 318 3400 430
rect 3350 272 3352 318
rect 3398 272 3400 318
rect 3350 210 3400 272
rect 3520 318 3570 380
rect 3520 272 3522 318
rect 3568 272 3570 318
rect 3520 140 3570 272
rect 3690 318 3740 970
rect 3690 272 3692 318
rect 3738 272 3740 318
rect 3690 210 3740 272
rect 0 118 3850 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1032 118
rect 1078 72 1262 118
rect 1308 72 1492 118
rect 1538 72 1722 118
rect 1768 72 1952 118
rect 1998 72 2182 118
rect 2228 72 2412 118
rect 2458 72 2642 118
rect 2688 72 2872 118
rect 2918 72 3102 118
rect 3148 72 3332 118
rect 3378 72 3562 118
rect 3608 72 3850 118
rect 0 0 3850 72
<< via1 >>
rect 134 992 142 1036
rect 142 992 186 1036
rect 134 984 186 992
rect 1374 854 1426 906
rect 554 773 606 776
rect 554 727 557 773
rect 557 727 603 773
rect 603 727 606 773
rect 554 724 606 727
rect 1104 773 1156 776
rect 1104 727 1107 773
rect 1107 727 1153 773
rect 1153 727 1156 773
rect 1104 724 1156 727
rect 2064 984 2116 1036
rect 1934 903 1986 906
rect 1934 857 1937 903
rect 1937 857 1983 903
rect 1983 857 1986 903
rect 1934 854 1986 857
rect 284 464 336 516
rect 794 464 846 516
rect 1534 513 1586 516
rect 1534 467 1537 513
rect 1537 467 1583 513
rect 1583 467 1586 513
rect 1534 464 1586 467
rect 2254 903 2306 906
rect 2254 857 2257 903
rect 2257 857 2303 903
rect 2303 857 2306 903
rect 2254 854 2306 857
rect 2834 984 2886 1036
rect 3204 984 3256 1036
rect 2504 854 2556 906
rect 2074 773 2126 776
rect 2074 727 2077 773
rect 2077 727 2123 773
rect 2123 727 2126 773
rect 2074 724 2126 727
rect 1934 643 1986 646
rect 1934 597 1937 643
rect 1937 597 1983 643
rect 1983 597 1986 643
rect 1934 594 1986 597
rect 2324 594 2376 646
rect 1874 334 1926 386
rect 3714 984 3766 1036
rect 3564 903 3616 906
rect 3564 857 3567 903
rect 3567 857 3613 903
rect 3613 857 3616 903
rect 3564 854 3616 857
rect 2654 602 2698 646
rect 2698 602 2706 646
rect 2654 594 2706 602
rect 3414 643 3466 646
rect 3414 597 3417 643
rect 3417 597 3463 643
rect 3463 597 3466 643
rect 3414 594 3466 597
rect 2834 503 2886 506
rect 2834 457 2837 503
rect 2837 457 2883 503
rect 2883 457 2886 503
rect 2834 454 2886 457
rect 3124 503 3176 506
rect 3124 457 3127 503
rect 3127 457 3173 503
rect 3173 457 3176 503
rect 3124 454 3176 457
<< metal2 >>
rect 110 1036 210 1050
rect 2050 1040 2130 1050
rect 2820 1040 2900 1050
rect 110 984 134 1036
rect 186 984 210 1036
rect 110 970 210 984
rect 2040 1036 2910 1040
rect 2040 984 2064 1036
rect 2116 984 2834 1036
rect 2886 984 2910 1036
rect 2040 980 2910 984
rect 3180 1036 3280 1050
rect 3700 1040 3780 1050
rect 3180 984 3204 1036
rect 3256 984 3280 1036
rect 2050 970 2130 980
rect 2820 970 2900 980
rect 3180 970 3280 984
rect 3690 1036 3790 1040
rect 3690 984 3714 1036
rect 3766 984 3790 1036
rect 3690 980 3790 984
rect 3700 970 3780 980
rect 1350 910 1440 920
rect 1910 910 2010 920
rect 2240 910 2320 920
rect 2490 910 2580 920
rect 3550 910 3630 920
rect 1350 906 2580 910
rect 1350 854 1374 906
rect 1426 854 1934 906
rect 1986 854 2254 906
rect 2306 854 2504 906
rect 2556 854 2580 906
rect 1350 850 2580 854
rect 3540 906 3640 910
rect 3540 854 3564 906
rect 3616 854 3640 906
rect 3540 850 3640 854
rect 1350 840 1440 850
rect 1910 840 2010 850
rect 2240 840 2320 850
rect 2490 840 2580 850
rect 3550 840 3630 850
rect 530 776 630 790
rect 530 724 554 776
rect 606 724 630 776
rect 530 710 630 724
rect 1080 776 1180 790
rect 2060 780 2140 790
rect 1080 724 1104 776
rect 1156 724 1180 776
rect 1080 710 1180 724
rect 2050 776 2150 780
rect 2050 724 2074 776
rect 2126 724 2150 776
rect 2050 720 2150 724
rect 2060 710 2140 720
rect 260 520 360 530
rect 550 520 610 710
rect 1920 650 2000 660
rect 2310 650 2390 660
rect 1910 646 2410 650
rect 1910 594 1934 646
rect 1986 594 2324 646
rect 2376 594 2410 646
rect 1910 590 2410 594
rect 2630 646 2730 660
rect 3400 650 3480 660
rect 2630 594 2654 646
rect 2706 594 2730 646
rect 1920 580 2000 590
rect 2310 580 2390 590
rect 2630 580 2730 594
rect 3330 646 3490 650
rect 3330 594 3414 646
rect 3466 594 3490 646
rect 3330 590 3490 594
rect 3400 580 3480 590
rect 260 516 610 520
rect 260 464 284 516
rect 336 464 610 516
rect 260 460 610 464
rect 260 450 360 460
rect 550 260 610 460
rect 770 520 870 530
rect 1520 520 1600 530
rect 770 516 1610 520
rect 770 464 794 516
rect 846 464 1534 516
rect 1586 464 1610 516
rect 770 460 1610 464
rect 2810 506 2910 520
rect 770 450 870 460
rect 1520 450 1600 460
rect 2810 454 2834 506
rect 2886 454 2910 506
rect 2810 440 2910 454
rect 3080 506 3200 520
rect 3080 454 3124 506
rect 3176 454 3200 506
rect 3080 440 3200 454
rect 1860 390 1940 400
rect 2810 390 2890 440
rect 1850 386 2890 390
rect 1850 334 1874 386
rect 1926 334 2890 386
rect 1850 330 2890 334
rect 1860 320 1940 330
rect 3080 260 3140 440
rect 550 200 3140 260
<< labels >>
rlabel via1 s 1104 724 1156 776 4 D
port 1 nsew signal input
rlabel via1 s 3714 984 3766 1036 4 Q
port 2 nsew signal output
rlabel via1 s 3564 854 3616 906 4 QN
port 3 nsew signal output
rlabel via1 s 134 984 186 1036 4 RN
port 4 nsew signal input
rlabel via1 s 2654 594 2706 646 4 CLK
port 5 nsew clock input
rlabel metal1 s 110 1110 160 1660 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 710 1110 760 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 980 1110 1030 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1590 1110 1640 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 1260 2200 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2680 1110 2730 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2920 1110 2970 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3520 1110 3570 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3850 1660 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 460 0 510 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 800 0 850 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 980 0 1030 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1590 0 1640 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2150 0 2200 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2680 0 2730 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2830 0 2880 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3170 0 3220 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3520 0 3570 380 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3850 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal2 s 2630 580 2730 660 1 CLK
port 5 nsew clock input
rlabel metal1 s 2630 590 2730 650 1 CLK
port 5 nsew clock input
rlabel metal2 s 1080 710 1180 790 1 D
port 1 nsew signal input
rlabel metal1 s 1080 720 1180 780 1 D
port 1 nsew signal input
rlabel metal2 s 3700 970 3780 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3690 980 3790 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 3690 210 3740 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 3690 970 3780 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 3690 980 3790 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 3550 840 3630 920 1 QN
port 3 nsew signal output
rlabel metal2 s 3540 850 3640 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3350 210 3400 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3350 850 3400 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 3350 430 3620 480 1 QN
port 3 nsew signal output
rlabel metal1 s 3570 430 3620 910 1 QN
port 3 nsew signal output
rlabel metal1 s 3350 850 3640 910 1 QN
port 3 nsew signal output
rlabel metal2 s 110 970 210 1050 1 RN
port 4 nsew signal input
rlabel metal1 s 110 980 210 1040 1 RN
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 3850 1660
string GDS_END 266902
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 239042
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
