VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__cor
  CLASS ENDCAP BOTTOMLEFT ;
  FOREIGN gf180mcu_fd_io__cor ;
  ORIGIN 0.000 0.000 ;
  SIZE 355.000 BY 355.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_COR_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 334.000 342.775 341.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.000 323.930 301.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 278.000 342.640 285.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 270.000 342.640 277.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262.000 342.640 269.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 214.000 342.640 229.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 290.485 214.000 353.065 228.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206.000 342.640 213.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 182.000 342.640 197.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 166.000 342.640 181.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 150.000 342.640 165.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 134.000 342.640 149.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.000 342.640 125.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 353.345 118.000 355.000 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 342.000 344.850 348.390 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.915 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 326.000 344.850 333.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.815 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 302.000 344.850 309.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.715 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.000 349.785 293.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 351.755 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 230.000 349.785 245.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.305 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 198.000 349.785 205.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 283.790 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126.000 349.785 133.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 253.700 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 102.000 349.785 117.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.045 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 86.000 349.785 101.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 269.350 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 349.785 85.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.045 70.000 355.000 85.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 310.000 352.150 317.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 342.635 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.000 307.295 261.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 342.635 254.000 355.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 65.540 65.540 355.000 355.000 ;
      LAYER Metal2 ;
        RECT 67.970 67.970 354.445 354.450 ;
      LAYER Metal3 ;
        RECT 246.800 347.985 252.200 352.200 ;
        RECT 318.800 350.350 324.200 352.200 ;
        RECT 70.000 340.840 116.200 347.985 ;
        RECT 126.800 340.840 132.200 347.985 ;
        RECT 198.800 340.840 204.200 347.985 ;
        RECT 230.800 340.840 252.200 347.985 ;
        RECT 286.800 340.840 292.200 347.985 ;
        RECT 310.800 343.050 324.200 350.350 ;
        RECT 350.190 350.190 355.000 354.000 ;
        RECT 70.000 305.495 252.200 340.840 ;
        RECT 262.800 322.130 292.200 340.840 ;
        RECT 302.800 340.975 332.200 343.050 ;
        RECT 342.800 340.975 350.115 343.050 ;
        RECT 302.800 340.200 350.115 340.975 ;
        RECT 302.800 334.800 351.545 340.200 ;
        RECT 302.800 324.200 350.015 334.800 ;
        RECT 302.800 322.130 352.200 324.200 ;
        RECT 262.800 318.800 352.200 322.130 ;
        RECT 262.800 308.200 340.835 318.800 ;
        RECT 262.800 305.495 349.915 308.200 ;
        RECT 70.000 300.200 349.915 305.495 ;
        RECT 70.000 294.800 351.545 300.200 ;
        RECT 70.000 284.200 349.955 294.800 ;
        RECT 70.000 262.800 351.545 284.200 ;
        RECT 70.000 252.200 340.835 262.800 ;
        RECT 70.000 246.800 352.200 252.200 ;
        RECT 70.000 230.795 295.505 246.800 ;
        RECT 70.000 212.200 288.685 230.795 ;
        RECT 354.865 214.800 355.000 228.200 ;
        RECT 70.000 206.800 351.545 212.200 ;
        RECT 70.000 196.200 281.990 206.800 ;
        RECT 70.000 134.800 351.545 196.200 ;
        RECT 70.000 124.200 251.900 134.800 ;
        RECT 70.000 118.800 351.545 124.200 ;
        RECT 70.000 102.800 284.245 118.800 ;
        RECT 70.000 84.200 267.550 102.800 ;
        RECT 70.000 70.000 284.245 84.200 ;
  END
END gf180mcu_fd_io__cor
END LIBRARY

