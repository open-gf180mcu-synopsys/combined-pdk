magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 1206 870
<< pwell >>
rect -86 -86 1206 352
<< mvnmos >>
rect 124 136 244 232
rect 348 136 468 232
rect 572 136 692 232
rect 796 136 916 232
<< mvpmos >>
rect 124 472 224 716
rect 368 472 468 716
rect 572 472 672 716
rect 816 472 916 716
<< mvndiff >>
rect 36 197 124 232
rect 36 151 49 197
rect 95 151 124 197
rect 36 136 124 151
rect 244 197 348 232
rect 244 151 273 197
rect 319 151 348 197
rect 244 136 348 151
rect 468 197 572 232
rect 468 151 497 197
rect 543 151 572 197
rect 468 136 572 151
rect 692 197 796 232
rect 692 151 721 197
rect 767 151 796 197
rect 692 136 796 151
rect 916 197 1004 232
rect 916 151 945 197
rect 991 151 1004 197
rect 916 136 1004 151
<< mvpdiff >>
rect 36 669 124 716
rect 36 529 49 669
rect 95 529 124 669
rect 36 472 124 529
rect 224 643 368 716
rect 224 503 273 643
rect 319 503 368 643
rect 224 472 368 503
rect 468 639 572 716
rect 468 593 497 639
rect 543 593 572 639
rect 468 472 572 593
rect 672 643 816 716
rect 672 503 721 643
rect 767 503 816 643
rect 672 472 816 503
rect 916 669 1004 716
rect 916 529 945 669
rect 991 529 1004 669
rect 916 472 1004 529
<< mvndiffc >>
rect 49 151 95 197
rect 273 151 319 197
rect 497 151 543 197
rect 721 151 767 197
rect 945 151 991 197
<< mvpdiffc >>
rect 49 529 95 669
rect 273 503 319 643
rect 497 593 543 639
rect 721 503 767 643
rect 945 529 991 669
<< polysilicon >>
rect 124 716 224 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 124 412 224 472
rect 368 412 468 472
rect 572 412 672 472
rect 816 412 916 472
rect 124 399 916 412
rect 124 353 203 399
rect 531 353 916 399
rect 124 335 916 353
rect 124 232 244 335
rect 348 232 468 335
rect 572 232 692 335
rect 796 232 916 335
rect 124 92 244 136
rect 348 92 468 136
rect 572 92 692 136
rect 796 92 916 136
<< polycontact >>
rect 203 353 531 399
<< metal1 >>
rect 0 724 1120 844
rect 49 669 95 724
rect 49 518 95 529
rect 273 643 319 654
rect 486 639 554 724
rect 945 669 991 724
rect 486 593 497 639
rect 543 593 554 639
rect 690 643 767 654
rect 690 541 721 643
rect 319 503 721 541
rect 945 518 991 529
rect 273 477 767 503
rect 130 399 542 430
rect 130 353 203 399
rect 531 353 542 399
rect 690 307 767 477
rect 273 243 767 307
rect 49 197 95 208
rect 49 60 95 151
rect 273 197 319 243
rect 690 197 767 243
rect 273 140 319 151
rect 486 151 497 197
rect 543 151 554 197
rect 486 60 554 151
rect 690 151 721 197
rect 690 140 767 151
rect 945 197 991 208
rect 945 60 991 151
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 600 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 945 197 991 208 0 FreeSans 600 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 690 541 767 654 0 FreeSans 600 0 0 0 ZN
port 2 nsew default output
flabel metal1 s 130 353 542 430 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 273 541 319 654 1 ZN
port 2 nsew default output
rlabel metal1 s 273 477 767 541 1 ZN
port 2 nsew default output
rlabel metal1 s 690 307 767 477 1 ZN
port 2 nsew default output
rlabel metal1 s 273 243 767 307 1 ZN
port 2 nsew default output
rlabel metal1 s 690 140 767 243 1 ZN
port 2 nsew default output
rlabel metal1 s 273 140 319 243 1 ZN
port 2 nsew default output
rlabel metal1 s 945 593 991 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 486 593 554 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 593 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 945 518 991 593 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 518 95 593 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 197 95 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1120 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string GDS_END 826338
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 823102
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
