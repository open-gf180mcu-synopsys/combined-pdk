magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_0
timestamp 1750858719
transform 1 0 11558 0 1 238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_1
timestamp 1750858719
transform 1 0 11558 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_2
timestamp 1750858719
transform 1 0 11558 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_3
timestamp 1750858719
transform 1 0 11935 0 1 22931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_4
timestamp 1750858719
transform 1 0 11935 0 1 23869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_5
timestamp 1750858719
transform 1 0 11935 0 1 24731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_6
timestamp 1750858719
transform 1 0 11935 0 1 25669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_7
timestamp 1750858719
transform 1 0 11935 0 1 26531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_8
timestamp 1750858719
transform 1 0 12313 0 1 21131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_9
timestamp 1750858719
transform 1 0 11935 0 1 28331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_10
timestamp 1750858719
transform 1 0 11935 0 1 27469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_11
timestamp 1750858719
transform 1 0 12691 0 1 7669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_12
timestamp 1750858719
transform 1 0 12691 0 1 8531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_13
timestamp 1750858719
transform 1 0 12691 0 1 9469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_14
timestamp 1750858719
transform 1 0 12691 0 1 10331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_15
timestamp 1750858719
transform 1 0 12691 0 1 11269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_16
timestamp 1750858719
transform 1 0 12691 0 1 12131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_17
timestamp 1750858719
transform 1 0 11558 0 1 28562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_18
timestamp 1750858719
transform 1 0 11558 0 1 26762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_19
timestamp 1750858719
transform 1 0 11558 0 1 24962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_20
timestamp 1750858719
transform 1 0 11558 0 1 23162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_21
timestamp 1750858719
transform 1 0 11558 0 1 21362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_22
timestamp 1750858719
transform 1 0 11558 0 1 19562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_23
timestamp 1750858719
transform 1 0 11558 0 1 17762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_24
timestamp 1750858719
transform 1 0 11558 0 1 15962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_25
timestamp 1750858719
transform 1 0 11558 0 1 14162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_26
timestamp 1750858719
transform 1 0 11558 0 1 12362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_27
timestamp 1750858719
transform 1 0 11558 0 1 10562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_28
timestamp 1750858719
transform 1 0 11558 0 1 8762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_29
timestamp 1750858719
transform 1 0 11558 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_30
timestamp 1750858719
transform 1 0 11558 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_31
timestamp 1750858719
transform 1 0 11558 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_32
timestamp 1750858719
transform 1 0 12313 0 1 14869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_33
timestamp 1750858719
transform 1 0 12313 0 1 15731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_34
timestamp 1750858719
transform 1 0 13068 0 1 6731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_35
timestamp 1750858719
transform 1 0 12313 0 1 16669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_36
timestamp 1750858719
transform 1 0 12691 0 1 13931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_37
timestamp 1750858719
transform 1 0 12691 0 1 13069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_38
timestamp 1750858719
transform 1 0 12313 0 1 17531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_39
timestamp 1750858719
transform 1 0 12313 0 1 18469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_40
timestamp 1750858719
transform 1 0 12313 0 1 19331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_41
timestamp 1750858719
transform 1 0 13068 0 1 469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_42
timestamp 1750858719
transform 1 0 13068 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_43
timestamp 1750858719
transform 1 0 13068 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_44
timestamp 1750858719
transform 1 0 13068 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_45
timestamp 1750858719
transform 1 0 13068 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_46
timestamp 1750858719
transform 1 0 13068 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_47
timestamp 1750858719
transform 1 0 13068 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_48
timestamp 1750858719
transform 1 0 11558 0 1 27238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_49
timestamp 1750858719
transform 1 0 11558 0 1 25438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_50
timestamp 1750858719
transform 1 0 11558 0 1 23638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_51
timestamp 1750858719
transform 1 0 11558 0 1 21838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_52
timestamp 1750858719
transform 1 0 11558 0 1 20038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_53
timestamp 1750858719
transform 1 0 11558 0 1 18238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_54
timestamp 1750858719
transform 1 0 11558 0 1 16438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_55
timestamp 1750858719
transform 1 0 11558 0 1 14638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_56
timestamp 1750858719
transform 1 0 11558 0 1 12838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_57
timestamp 1750858719
transform 1 0 11558 0 1 11038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_58
timestamp 1750858719
transform 1 0 11558 0 1 9238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_59
timestamp 1750858719
transform 1 0 11558 0 1 7438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_60
timestamp 1750858719
transform 1 0 11558 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_61
timestamp 1750858719
transform 1 0 11558 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_62
timestamp 1750858719
transform 1 0 12313 0 1 20269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_63
timestamp 1750858719
transform 1 0 11935 0 1 22069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_64
timestamp 1750858719
transform 1 0 17864 0 1 578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_65
timestamp 1750858719
transform 1 0 17487 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_66
timestamp 1750858719
transform 1 0 17109 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_67
timestamp 1750858719
transform 1 0 16731 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_68
timestamp 1750858719
transform 1 0 16354 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_69
timestamp 1750858719
transform 1 0 15976 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_70
timestamp 1750858719
transform 1 0 15598 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_71
timestamp 1750858719
transform 1 0 15220 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_72
timestamp 1750858719
transform 1 0 15220 0 1 13822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_73
timestamp 1750858719
transform 1 0 15220 0 1 21022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_74
timestamp 1750858719
transform 1 0 15220 0 1 28222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_75
timestamp 1750858719
transform 1 0 15598 0 1 13178
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_76
timestamp 1750858719
transform 1 0 15598 0 1 20378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_77
timestamp 1750858719
transform 1 0 15598 0 1 27578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_78
timestamp 1750858719
transform 1 0 15976 0 1 12022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_79
timestamp 1750858719
transform 1 0 15976 0 1 19222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_80
timestamp 1750858719
transform 1 0 15976 0 1 26422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_81
timestamp 1750858719
transform 1 0 16354 0 1 11378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_82
timestamp 1750858719
transform 1 0 16354 0 1 18578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_83
timestamp 1750858719
transform 1 0 16354 0 1 25778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_84
timestamp 1750858719
transform 1 0 16731 0 1 10222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_85
timestamp 1750858719
transform 1 0 16731 0 1 17422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_86
timestamp 1750858719
transform 1 0 16731 0 1 24622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_87
timestamp 1750858719
transform 1 0 17109 0 1 9578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_88
timestamp 1750858719
transform 1 0 17109 0 1 16778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_89
timestamp 1750858719
transform 1 0 17109 0 1 23978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_90
timestamp 1750858719
transform 1 0 17487 0 1 8422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_91
timestamp 1750858719
transform 1 0 17487 0 1 15622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_92
timestamp 1750858719
transform 1 0 17487 0 1 22822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_93
timestamp 1750858719
transform 1 0 17864 0 1 7778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_94
timestamp 1750858719
transform 1 0 17864 0 1 14978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_95
timestamp 1750858719
transform 1 0 17864 0 1 22178
box 0 0 1 1
use xdec8_512x8m81  xdec8_512x8m81_0
timestamp 1750858719
transform 1 0 0 0 1 21600
box 1426 -1 22889 7201
use xdec8_512x8m81  xdec8_512x8m81_1
timestamp 1750858719
transform 1 0 0 0 1 0
box 1426 -1 22889 7201
use xdec8_512x8m81  xdec8_512x8m81_2
timestamp 1750858719
transform 1 0 0 0 1 7200
box 1426 -1 22889 7201
use xdec8_512x8m81  xdec8_512x8m81_3
timestamp 1750858719
transform 1 0 0 0 1 14400
box 1426 -1 22889 7201
<< properties >>
string GDS_END 2447752
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2434302
<< end >>
