magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< metal1 >>
rect 282 67176 86090 67894
rect 282 1000 1000 67176
rect 85372 1000 86090 67176
rect 282 282 86090 1000
<< obsm1 >>
rect 1000 1000 85372 67176
<< metal2 >>
rect 282 67568 86090 67894
rect 706 67176 86090 67376
rect 282 65478 606 66174
rect 282 63678 606 64374
rect 282 61878 606 62574
rect 282 60078 606 60774
rect 282 58278 606 58974
rect 282 56478 606 57174
rect 282 54678 606 55374
rect 282 52878 606 53574
rect 282 51078 606 51774
rect 282 49278 606 49974
rect 282 47478 606 48174
rect 282 45678 606 46374
rect 282 43878 606 44574
rect 282 42078 606 42774
rect 282 40278 606 40974
rect 282 38478 606 39174
rect 282 36678 606 37374
rect 282 34578 606 35274
rect 282 26538 606 28350
rect 282 21311 606 22255
rect 282 14398 606 17698
rect 282 10227 606 11419
rect 282 5771 606 7583
rect 282 2527 606 3719
rect 706 1000 1000 67176
rect 85372 66376 86090 67176
rect 85372 1000 85666 66376
rect 85766 65478 86090 66174
rect 85766 63678 86090 64374
rect 85766 61878 86090 62574
rect 85766 60078 86090 60774
rect 85766 58278 86090 58974
rect 85766 56478 86090 57174
rect 85766 54678 86090 55374
rect 85766 52878 86090 53574
rect 85766 51078 86090 51774
rect 85766 49278 86090 49974
rect 85766 47478 86090 48174
rect 85766 45678 86090 46374
rect 85766 43878 86090 44574
rect 85766 42078 86090 42774
rect 85766 40278 86090 40974
rect 85766 38478 86090 39174
rect 85766 36678 86090 37374
rect 85766 34578 86090 35274
rect 85766 26538 86090 28350
rect 85766 21311 86090 22255
rect 85766 14398 86090 17698
rect 85766 10227 86090 11419
rect 85766 5771 86090 7583
rect 85766 2527 86090 3719
rect 706 282 1706 1000
rect 1864 0 2088 1000
rect 2539 0 2763 1000
rect 3380 0 3604 1000
rect 4642 282 5642 1000
rect 6927 282 7151 1000
rect 7946 282 8170 1000
rect 9442 282 10442 1000
rect 11533 0 11757 1000
rect 12206 0 12430 1000
rect 12604 0 12828 1000
rect 13054 0 13278 1000
rect 13454 0 13678 1000
rect 14127 0 14351 1000
rect 15442 282 16442 1000
rect 17727 282 17951 1000
rect 18746 282 18970 1000
rect 20242 282 21242 1000
rect 22279 0 22503 1000
rect 23404 0 23628 1000
rect 23795 0 24019 1000
rect 24856 282 25080 1000
rect 25873 282 26097 1000
rect 27936 0 28160 1000
rect 29006 0 29230 1000
rect 29705 0 29929 1000
rect 30859 0 31083 1000
rect 31324 282 32324 1000
rect 32552 0 32776 1000
rect 33022 282 34022 1000
rect 34243 0 34467 1000
rect 34831 282 35831 1000
rect 38028 282 39028 1000
rect 40588 0 40812 1000
rect 41233 282 42233 1000
rect 43633 282 44633 1000
rect 46033 282 47033 1000
rect 50342 0 50566 1000
rect 51233 282 52233 1000
rect 52478 282 53478 1000
rect 53772 0 53996 1000
rect 54417 0 54641 1000
rect 55164 0 55388 1000
rect 56265 0 56489 1000
rect 59313 282 59537 1000
rect 60330 282 60554 1000
rect 61447 0 61671 1000
rect 62115 0 62339 1000
rect 62958 0 63182 1000
rect 64218 282 65218 1000
rect 66502 282 66726 1000
rect 67521 282 67745 1000
rect 69018 282 70018 1000
rect 71109 0 71333 1000
rect 71782 0 72006 1000
rect 72180 0 72404 1000
rect 72630 0 72854 1000
rect 73030 0 73254 1000
rect 73703 0 73927 1000
rect 75018 282 76018 1000
rect 77301 282 77525 1000
rect 78320 282 78544 1000
rect 79818 282 80818 1000
rect 81855 0 82079 1000
rect 82695 0 82919 1000
rect 83372 0 83596 1000
rect 84666 282 85666 1000
<< obsm2 >>
rect 1000 1000 85372 67176
<< metal3 >>
rect 1401 67376 2401 68176
rect 2626 67568 3626 68176
rect 4137 67376 5137 68176
rect 5362 67568 6362 68176
rect 6801 67376 7801 68176
rect 8026 67568 9026 68176
rect 9537 67376 10537 68176
rect 10762 67568 11762 68176
rect 12201 67376 13201 68176
rect 13426 67568 14426 68176
rect 14937 67376 15937 68176
rect 16162 67568 17162 68176
rect 17601 67376 18601 68176
rect 18826 67568 19826 68176
rect 20653 67376 21653 68176
rect 22258 67568 23258 68176
rect 23483 67376 24483 68176
rect 25158 67568 26158 68176
rect 26572 67376 27572 68176
rect 27877 67568 28877 68176
rect 29273 67568 30273 68176
rect 30710 67376 31710 68176
rect 32381 67568 33381 68176
rect 34024 67568 35024 68176
rect 35415 67376 36415 68176
rect 36948 67568 37948 68176
rect 38585 67376 39585 68176
rect 39882 67568 40882 68176
rect 41230 67376 42230 68176
rect 42430 67568 43430 68176
rect 43713 67568 44713 68176
rect 45069 67376 46069 68176
rect 46313 67376 47313 68176
rect 47538 67568 48538 68176
rect 48901 67376 49901 68176
rect 50465 67568 51465 68176
rect 52569 67376 53569 68176
rect 54262 67376 55262 68176
rect 55990 67568 56990 68176
rect 57547 67376 58547 68176
rect 58791 67568 59791 68176
rect 60977 67376 61977 68176
rect 62202 67568 63202 68176
rect 63713 67376 64713 68176
rect 64938 67568 65938 68176
rect 66377 67568 67378 68176
rect 67602 67568 68603 68176
rect 66378 67376 67378 67568
rect 69113 67376 70113 68176
rect 70338 67568 71338 68176
rect 71777 67376 72777 68176
rect 73002 67568 74002 68176
rect 74513 67376 75513 68176
rect 75738 67568 76738 68176
rect 77177 67376 78177 68176
rect 78402 67568 79402 68176
rect 80229 67376 81229 68176
rect 81834 67568 82834 68176
rect 83059 67376 84059 68176
rect 84666 67376 85666 68176
rect 0 67176 86372 67376
rect 0 66376 1000 67176
rect 0 65476 1000 66176
rect 85372 66376 86372 67176
rect 30402 65726 54622 65928
rect 85372 65476 86372 66176
rect 0 64576 1706 65276
rect 85372 64576 86372 65276
rect 0 63676 1000 64376
rect 30403 63926 54622 64128
rect 0 62776 1000 63476
rect 0 61876 1000 62576
rect 85372 63676 86372 64376
rect 85372 62776 86372 63476
rect 30403 62126 54622 62328
rect 0 60976 1000 61676
rect 0 60076 1000 60776
rect 85372 61876 86372 62576
rect 85372 60976 86372 61676
rect 30403 60326 54622 60528
rect 0 59176 1000 59876
rect 0 58276 1000 58976
rect 85372 60076 86372 60776
rect 85372 59176 86372 59876
rect 30403 58526 54622 58728
rect 0 57376 1000 58076
rect 0 56476 1000 57176
rect 85372 58276 86372 58976
rect 85372 57376 86372 58076
rect 30403 56726 54622 56928
rect 0 55576 1000 56276
rect 0 54676 1000 55376
rect 85372 56476 86372 57176
rect 85372 55576 86372 56276
rect 30403 54926 54622 55128
rect 0 53776 1000 54476
rect 0 52876 1000 53576
rect 85372 54676 86372 55376
rect 85372 53776 86372 54476
rect 30403 53126 54622 53328
rect 0 51976 1000 52676
rect 0 51076 1000 51776
rect 85372 52876 86372 53576
rect 85372 51976 86372 52676
rect 30403 51326 54622 51528
rect 0 50176 1000 50876
rect 0 49276 1000 49976
rect 85372 51076 86372 51776
rect 85372 50176 86372 50876
rect 30403 49526 54622 49728
rect 0 48376 1000 49076
rect 0 47476 1000 48176
rect 85372 49276 86372 49976
rect 85372 48376 86372 49076
rect 30403 47726 54622 47928
rect 0 46576 1000 47276
rect 0 45676 1000 46376
rect 85372 47476 86372 48176
rect 85372 46576 86372 47276
rect 30403 45926 54622 46128
rect 0 44776 1000 45476
rect 0 43876 1000 44576
rect 85372 45676 86372 46376
rect 85372 44776 86372 45476
rect 30403 44126 54622 44328
rect 0 42976 1000 43676
rect 0 42076 1000 42776
rect 85372 43876 86372 44576
rect 85372 42976 86372 43676
rect 30403 42326 54622 42528
rect 0 41176 1000 41876
rect 0 40276 1000 40976
rect 85372 42076 86372 42776
rect 85372 41176 86372 41876
rect 30403 40526 54622 40728
rect 0 39376 1000 40076
rect 0 38476 1000 39176
rect 85372 40276 86372 40976
rect 85372 39376 86372 40076
rect 30403 38726 54622 38928
rect 0 37576 1000 38276
rect 0 36676 1000 37376
rect 85372 38476 86372 39176
rect 85372 37576 86372 38276
rect 30403 36926 54622 37128
rect 0 35776 1000 36476
rect 85372 36676 86372 37376
rect 85372 35776 86372 36476
rect 0 34536 1000 35326
rect 27442 34494 27782 35062
rect 60559 34536 60647 35387
rect 85372 34536 86372 35326
rect 0 29430 1000 34125
rect 2095 32315 2188 34126
rect 61853 32315 72383 34125
rect 26772 31486 58351 32199
rect 0 26435 1000 28416
rect 1954 26435 26070 28434
rect 26772 27382 58351 30105
rect 85372 29430 86372 34125
rect 58785 26435 84717 28434
rect 85372 26435 86372 28416
rect 0 22938 1000 23938
rect 26770 23370 58348 24278
rect 0 21282 1000 22282
rect 24036 21826 27826 22282
rect 56078 21826 57677 23199
rect 85372 22938 86372 23938
rect 0 18016 1000 20739
rect 29513 19969 55645 21625
rect 85372 21282 86372 22282
rect 61502 18015 83763 20739
rect 85372 18016 86372 20739
rect 0 14328 1000 17730
rect 24111 14329 27828 16598
rect 0 12036 1000 14178
rect 29478 13243 45977 15015
rect 57295 14327 83763 16784
rect 85372 14328 86372 17730
rect 23821 12046 34761 12847
rect 50228 12035 58421 13866
rect 59826 12035 60026 14017
rect 61807 13461 72429 14178
rect 83169 13461 84221 14179
rect 83169 12035 84221 12847
rect 85372 12036 86372 14178
rect 0 10176 1000 11493
rect 2249 10174 24250 11491
rect 42261 10740 57736 11527
rect 0 8152 1000 9515
rect 2226 8154 28729 9515
rect 41857 9165 51430 10420
rect 60736 10173 84482 11491
rect 85372 10176 86372 11493
rect 29513 7900 41397 8582
rect 57909 8154 62278 9516
rect 72602 8152 83234 9515
rect 85372 8152 86372 9515
rect 0 5766 1000 7596
rect 2249 6980 24250 7595
rect 29537 6744 34622 7652
rect 34860 6592 55482 7392
rect 60736 6980 84787 7595
rect 23687 6177 41397 6199
rect 50922 5766 62429 6199
rect 85372 5766 86372 7596
rect 0 4060 1000 5629
rect 23687 5175 27214 5630
rect 57909 5175 62429 5630
rect 23909 4166 62429 4619
rect 85372 4060 86372 5629
rect 0 2502 1000 3772
rect 27438 3524 27778 3876
rect 28764 3524 28894 3876
rect 41774 3524 41904 3876
rect 42299 3524 42429 3876
rect 46873 3524 47003 3876
rect 47321 3524 47451 3876
rect 47769 3524 47899 3876
rect 48217 3524 48347 3876
rect 57345 3524 61215 3876
rect 0 1232 1000 2232
rect 706 1000 1000 1232
rect 85372 2502 86372 3772
rect 85372 1232 86372 2232
rect 85372 1000 85666 1232
rect 706 0 1706 1000
rect 2039 0 3039 1000
rect 3442 0 4442 1000
rect 4642 0 5642 932
rect 5842 0 6842 1000
rect 7042 0 8042 1000
rect 8242 0 9242 1000
rect 9442 0 10442 932
rect 10642 0 11642 1000
rect 12443 0 13443 1000
rect 14242 0 15242 1000
rect 15442 0 16442 932
rect 16642 0 17642 1000
rect 17842 0 18842 1000
rect 19042 0 20042 1000
rect 20242 0 21242 932
rect 21910 0 22910 1000
rect 23110 0 24110 1000
rect 24410 0 25410 1000
rect 25710 0 26710 1000
rect 27010 0 28010 1000
rect 28310 0 29310 1000
rect 29610 0 30610 1000
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1000
rect 38028 0 39028 932
rect 39228 0 40228 1000
rect 41233 0 42233 932
rect 42433 0 43433 1000
rect 43633 0 44633 932
rect 44833 0 45833 1000
rect 46033 0 47033 932
rect 47233 0 48233 1000
rect 48566 0 49566 1000
rect 49876 0 50876 1000
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1000
rect 55758 0 56758 1000
rect 57058 0 58058 1000
rect 58358 0 59358 1000
rect 59658 0 60658 1000
rect 60958 0 61958 1000
rect 62295 0 63295 1000
rect 64218 0 65218 932
rect 65418 0 66418 1000
rect 66618 0 67618 1000
rect 67818 0 68818 1000
rect 69018 0 70018 932
rect 70218 0 71218 1000
rect 72017 0 73017 1000
rect 73818 0 74818 1000
rect 75018 0 76018 932
rect 76218 0 77218 1000
rect 77418 0 78418 1000
rect 78618 0 79618 1000
rect 79818 0 80818 932
rect 81018 0 82018 1000
rect 82419 0 83419 1000
rect 84666 0 85666 1000
<< obsm3 >>
rect 1000 65928 85372 67176
rect 1000 65726 30402 65928
rect 54622 65726 85372 65928
rect 1000 65276 85372 65726
rect 1706 64576 85372 65276
rect 1000 64128 85372 64576
rect 1000 63926 30403 64128
rect 54622 63926 85372 64128
rect 1000 62328 85372 63926
rect 1000 62126 30403 62328
rect 54622 62126 85372 62328
rect 1000 60528 85372 62126
rect 1000 60326 30403 60528
rect 54622 60326 85372 60528
rect 1000 58728 85372 60326
rect 1000 58526 30403 58728
rect 54622 58526 85372 58728
rect 1000 56928 85372 58526
rect 1000 56726 30403 56928
rect 54622 56726 85372 56928
rect 1000 55128 85372 56726
rect 1000 54926 30403 55128
rect 54622 54926 85372 55128
rect 1000 53328 85372 54926
rect 1000 53126 30403 53328
rect 54622 53126 85372 53328
rect 1000 51528 85372 53126
rect 1000 51326 30403 51528
rect 54622 51326 85372 51528
rect 1000 49728 85372 51326
rect 1000 49526 30403 49728
rect 54622 49526 85372 49728
rect 1000 47928 85372 49526
rect 1000 47726 30403 47928
rect 54622 47726 85372 47928
rect 1000 46128 85372 47726
rect 1000 45926 30403 46128
rect 54622 45926 85372 46128
rect 1000 44328 85372 45926
rect 1000 44126 30403 44328
rect 54622 44126 85372 44328
rect 1000 42528 85372 44126
rect 1000 42326 30403 42528
rect 54622 42326 85372 42528
rect 1000 40728 85372 42326
rect 1000 40526 30403 40728
rect 54622 40526 85372 40728
rect 1000 38928 85372 40526
rect 1000 38726 30403 38928
rect 54622 38726 85372 38928
rect 1000 37128 85372 38726
rect 1000 36926 30403 37128
rect 54622 36926 85372 37128
rect 1000 35387 85372 36926
rect 1000 35062 60559 35387
rect 1000 34494 27442 35062
rect 27782 34536 60559 35062
rect 60647 34536 85372 35387
rect 27782 34494 85372 34536
rect 1000 34126 85372 34494
rect 1000 32315 2095 34126
rect 2188 34125 85372 34126
rect 2188 32315 61853 34125
rect 72383 32315 85372 34125
rect 1000 32199 85372 32315
rect 1000 31486 26772 32199
rect 58351 31486 85372 32199
rect 1000 30105 85372 31486
rect 1000 28434 26772 30105
rect 1000 26435 1954 28434
rect 26070 27382 26772 28434
rect 58351 28434 85372 30105
rect 58351 27382 58785 28434
rect 26070 26435 58785 27382
rect 84717 26435 85372 28434
rect 1000 24278 85372 26435
rect 1000 23370 26770 24278
rect 58348 23370 85372 24278
rect 1000 23199 85372 23370
rect 1000 22282 56078 23199
rect 1000 21826 24036 22282
rect 27826 21826 56078 22282
rect 57677 21826 85372 23199
rect 1000 21625 85372 21826
rect 1000 19969 29513 21625
rect 55645 20739 85372 21625
rect 55645 19969 61502 20739
rect 1000 18015 61502 19969
rect 83763 18015 85372 20739
rect 1000 16784 85372 18015
rect 1000 16598 57295 16784
rect 1000 14329 24111 16598
rect 27828 15015 57295 16598
rect 27828 14329 29478 15015
rect 1000 13243 29478 14329
rect 45977 14327 57295 15015
rect 83763 14327 85372 16784
rect 45977 14179 85372 14327
rect 45977 14178 83169 14179
rect 45977 14017 61807 14178
rect 45977 13866 59826 14017
rect 45977 13243 50228 13866
rect 1000 12847 50228 13243
rect 1000 12046 23821 12847
rect 34761 12046 50228 12847
rect 1000 12035 50228 12046
rect 58421 12035 59826 13866
rect 60026 13461 61807 14017
rect 72429 13461 83169 14178
rect 84221 13461 85372 14179
rect 60026 12847 85372 13461
rect 60026 12035 83169 12847
rect 84221 12035 85372 12847
rect 1000 11527 85372 12035
rect 1000 11491 42261 11527
rect 1000 10174 2249 11491
rect 24250 10740 42261 11491
rect 57736 11491 85372 11527
rect 57736 10740 60736 11491
rect 24250 10420 60736 10740
rect 24250 10174 41857 10420
rect 1000 9515 41857 10174
rect 1000 8154 2226 9515
rect 28729 9165 41857 9515
rect 51430 10173 60736 10420
rect 84482 10173 85372 11491
rect 51430 9516 85372 10173
rect 51430 9165 57909 9516
rect 28729 8582 57909 9165
rect 28729 8154 29513 8582
rect 1000 7900 29513 8154
rect 41397 8154 57909 8582
rect 62278 9515 85372 9516
rect 62278 8154 72602 9515
rect 41397 8152 72602 8154
rect 83234 8152 85372 9515
rect 41397 7900 85372 8152
rect 1000 7652 85372 7900
rect 1000 7595 29537 7652
rect 1000 6980 2249 7595
rect 24250 6980 29537 7595
rect 1000 6744 29537 6980
rect 34622 7595 85372 7652
rect 34622 7392 60736 7595
rect 34622 6744 34860 7392
rect 1000 6592 34860 6744
rect 55482 6980 60736 7392
rect 84787 6980 85372 7595
rect 55482 6592 85372 6980
rect 1000 6199 85372 6592
rect 1000 6177 23687 6199
rect 41397 6177 50922 6199
rect 1000 5766 50922 6177
rect 62429 5766 85372 6199
rect 1000 5630 85372 5766
rect 1000 5175 23687 5630
rect 27214 5175 57909 5630
rect 62429 5175 85372 5630
rect 1000 4619 85372 5175
rect 1000 4166 23909 4619
rect 62429 4166 85372 4619
rect 1000 3876 85372 4166
rect 1000 3524 27438 3876
rect 27778 3524 28764 3876
rect 28894 3524 41774 3876
rect 41904 3524 42299 3876
rect 42429 3524 46873 3876
rect 47003 3524 47321 3876
rect 47451 3524 47769 3876
rect 47899 3524 48217 3876
rect 48347 3524 57345 3876
rect 61215 3524 85372 3876
rect 1000 1000 85372 3524
<< labels >>
rlabel metal2 s 29705 0 29929 1000 6 A[7]
port 1 nsew signal input
rlabel metal2 s 53772 0 53996 1000 6 A[6]
port 2 nsew signal input
rlabel metal2 s 54417 0 54641 1000 6 A[5]
port 3 nsew signal input
rlabel metal2 s 55164 0 55388 1000 6 A[4]
port 4 nsew signal input
rlabel metal2 s 56265 0 56489 1000 6 A[3]
port 5 nsew signal input
rlabel metal2 s 30859 0 31083 1000 6 A[2]
port 6 nsew signal input
rlabel metal2 s 32552 0 32776 1000 6 A[1]
port 7 nsew signal input
rlabel metal2 s 34243 0 34467 1000 6 A[0]
port 8 nsew signal input
rlabel metal2 s 50342 0 50566 1000 6 CEN
port 9 nsew signal input
rlabel metal2 s 27936 0 28160 1000 6 CLK
port 10 nsew signal input
rlabel metal2 s 83372 0 83596 1000 6 D[7]
port 11 nsew signal input
rlabel metal2 s 73030 0 73254 1000 6 D[6]
port 12 nsew signal input
rlabel metal2 s 71782 0 72006 1000 6 D[5]
port 13 nsew signal input
rlabel metal2 s 61447 0 61671 1000 6 D[4]
port 14 nsew signal input
rlabel metal2 s 23795 0 24019 1000 6 D[3]
port 15 nsew signal input
rlabel metal2 s 13454 0 13678 1000 6 D[2]
port 16 nsew signal input
rlabel metal2 s 12206 0 12430 1000 6 D[1]
port 17 nsew signal input
rlabel metal2 s 1864 0 2088 1000 6 D[0]
port 18 nsew signal input
rlabel metal2 s 40588 0 40812 1000 6 GWEN
port 19 nsew signal input
rlabel metal2 s 81855 0 82079 1000 6 Q[7]
port 20 nsew signal output
rlabel metal2 s 73703 0 73927 1000 6 Q[6]
port 21 nsew signal output
rlabel metal2 s 71109 0 71333 1000 6 Q[5]
port 22 nsew signal output
rlabel metal2 s 62958 0 63182 1000 6 Q[4]
port 23 nsew signal output
rlabel metal2 s 22279 0 22503 1000 6 Q[3]
port 24 nsew signal output
rlabel metal2 s 14127 0 14351 1000 6 Q[2]
port 25 nsew signal output
rlabel metal2 s 11533 0 11757 1000 6 Q[1]
port 26 nsew signal output
rlabel metal2 s 3380 0 3604 1000 6 Q[0]
port 27 nsew signal output
rlabel metal3 s 84666 0 85666 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 82419 0 83419 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 81018 0 82018 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 78618 0 79618 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 77418 0 78418 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 76218 0 77218 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 73818 0 74818 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 72017 0 73017 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 70218 0 71218 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 67818 0 68818 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 66618 0 67618 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 65418 0 66418 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 62295 0 63295 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 60958 0 61958 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 59658 0 60658 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 58358 0 59358 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57058 0 58058 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 55758 0 56758 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 54458 0 55458 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 49876 0 50876 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 48566 0 49566 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 47233 0 48233 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 44833 0 45833 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 42433 0 43433 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 39228 0 40228 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 36031 0 37031 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 29610 0 30610 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 28310 0 29310 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 27010 0 28010 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 25710 0 26710 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 24410 0 25410 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23110 0 24110 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 21910 0 22910 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 19042 0 20042 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 17842 0 18842 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 16642 0 17642 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 14242 0 15242 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 12443 0 13443 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 10642 0 11642 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 8242 0 9242 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 7042 0 8042 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 5842 0 6842 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 3442 0 4442 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 2039 0 3039 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 706 0 1706 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 1000 85666 1232 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 1232 86372 2232 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 706 1000 1000 1232 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 1232 1000 2232 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 4060 86372 5629 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 4060 1000 5629 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 8152 86372 9515 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 8152 1000 9515 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 12036 86372 14178 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 12036 1000 14178 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 18016 86372 20739 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 18016 1000 20739 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 22938 86372 23938 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 22938 1000 23938 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 29430 86372 34125 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 29430 1000 34125 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 35776 86372 36476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 35776 1000 36476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 37576 86372 38276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 37576 1000 38276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 39376 86372 40076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 39376 1000 40076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 41176 86372 41876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 41176 1000 41876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 42976 86372 43676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 42976 1000 43676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 44776 86372 45476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 44776 1000 45476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 46576 86372 47276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 46576 1000 47276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 48376 86372 49076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 48376 1000 49076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 50176 86372 50876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 50176 1000 50876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 51976 86372 52676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 51976 1000 52676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 53776 86372 54476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 53776 1000 54476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 55576 86372 56276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 55576 1000 56276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 57376 86372 58076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 57376 1000 58076 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 59176 86372 59876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 59176 1000 59876 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 60976 86372 61676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 60976 1000 61676 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 62776 86372 63476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 62776 1000 63476 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 64576 86372 65276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 64576 1706 65276 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 85372 66376 86372 67176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 66376 1000 67176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 67176 86372 67376 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 84666 67376 85666 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 83059 67376 84059 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 80229 67376 81229 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 77177 67376 78177 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 74513 67376 75513 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 71777 67376 72777 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 69113 67376 70113 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 66378 67376 67378 67568 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 66377 67568 67378 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 63713 67376 64713 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 60977 67376 61977 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57547 67376 58547 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 54262 67376 55262 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 52569 67376 53569 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 48901 67376 49901 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 46313 67376 47313 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 45069 67376 46069 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 41230 67376 42230 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 38585 67376 39585 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 35415 67376 36415 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 30710 67376 31710 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 26572 67376 27572 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23483 67376 24483 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 20653 67376 21653 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 17601 67376 18601 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 14937 67376 15937 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 12201 67376 13201 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 9537 67376 10537 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 6801 67376 7801 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 4137 67376 5137 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 1401 67376 2401 68176 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 84666 282 85666 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 706 282 1706 1000 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 85372 1000 85666 66376 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 85372 66376 86090 67176 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 706 1000 1000 67176 6 VDD
port 28 nsew power bidirectional
rlabel metal2 s 706 67176 86090 67376 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 2226 8154 28729 9515 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 29537 6744 34622 7652 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 2095 32315 2188 34126 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 26772 31486 58351 32199 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 26772 27382 58351 30105 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 61853 32315 72383 34125 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 26770 23370 58348 24278 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 29513 19969 55645 21625 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 61502 18015 83763 20739 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23821 12046 34761 12847 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 50228 12035 58421 13866 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 59826 12035 60026 14017 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 61807 13461 72429 14178 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 83169 12035 84221 12847 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 83169 13461 84221 14179 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57909 8154 62278 9516 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 72602 8152 83234 9515 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 6 VDD
port 28 nsew power bidirectional
rlabel metal3 s 79818 0 80818 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 75018 0 76018 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 69018 0 70018 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 64218 0 65218 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 52478 0 53478 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 51233 0 52233 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 46033 0 47033 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 43633 0 44633 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41233 0 42233 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 38028 0 39028 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 34831 0 35831 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 33022 0 34022 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 31324 0 32324 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 20242 0 21242 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 15442 0 16442 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 9442 0 10442 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 4642 0 5642 932 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 2502 86372 3772 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 5766 86372 7596 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 5766 1000 7596 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 10176 86372 11493 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 10176 1000 11493 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 14328 86372 17730 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14328 1000 17730 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 21282 86372 22282 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 21282 1000 22282 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 26435 86372 28416 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 26435 1000 28416 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 34536 86372 35326 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 34536 1000 35326 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 36676 86372 37376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 36676 1000 37376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 38476 86372 39176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 38476 1000 39176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 40276 86372 40976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 40276 1000 40976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 42076 86372 42776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 42076 1000 42776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 43876 86372 44576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 43876 1000 44576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 45676 86372 46376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 45676 1000 46376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 47476 86372 48176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 47476 1000 48176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 49276 86372 49976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 49276 1000 49976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 51076 86372 51776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 51076 1000 51776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 52876 86372 53576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 52876 1000 53576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 54676 86372 55376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 54676 1000 55376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 56476 86372 57176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 56476 1000 57176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 58276 86372 58976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 58276 1000 58976 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 60076 86372 60776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 60076 1000 60776 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 61876 86372 62576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 61876 1000 62576 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 63676 86372 64376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 63676 1000 64376 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85372 65476 86372 66176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 65476 1000 66176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 81834 67568 82834 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 78402 67568 79402 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 75738 67568 76738 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 73002 67568 74002 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 70338 67568 71338 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 67602 67568 68603 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 64938 67568 65938 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 62202 67568 63202 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 58791 67568 59791 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 55990 67568 56990 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50465 67568 51465 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 47538 67568 48538 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 43713 67568 44713 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 42430 67568 43430 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 39882 67568 40882 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 36948 67568 37948 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 34024 67568 35024 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 32381 67568 33381 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29273 67568 30273 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27877 67568 28877 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 25158 67568 26158 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 22258 67568 23258 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 18826 67568 19826 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 16162 67568 17162 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 13426 67568 14426 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 10762 67568 11762 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 8026 67568 9026 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 5362 67568 6362 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 2626 67568 3626 68176 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 79818 282 80818 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 78320 282 78544 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 77301 282 77525 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 75018 282 76018 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 69018 282 70018 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 67521 282 67745 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 66502 282 66726 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 64218 282 65218 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 60330 282 60554 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 59313 282 59537 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 52478 282 53478 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 51233 282 52233 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 46033 282 47033 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 43633 282 44633 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 41233 282 42233 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 38028 282 39028 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 34831 282 35831 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 33022 282 34022 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 31324 282 32324 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 29006 0 29230 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 25873 282 26097 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 24856 282 25080 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 20242 282 21242 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 18746 282 18970 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 17727 282 17951 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 15442 282 16442 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 9442 282 10442 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 7946 282 8170 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 6927 282 7151 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 4642 282 5642 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 2527 86090 3719 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 2527 606 3719 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 5771 86090 7583 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 5771 606 7583 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 10227 86090 11419 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 10227 606 11419 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 14398 86090 17698 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 14398 606 17698 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 21311 86090 22255 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 21311 606 22255 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 26538 86090 28350 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 26538 606 28350 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 34578 86090 35274 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 34578 606 35274 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 36678 86090 37374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 36678 606 37374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 38478 86090 39174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 38478 606 39174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 40278 86090 40974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 40278 606 40974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 42078 86090 42774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 42078 606 42774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 43878 86090 44574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 43878 606 44574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 45678 86090 46374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 45678 606 46374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 47478 86090 48174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 47478 606 48174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 49278 86090 49974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 49278 606 49974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 51078 86090 51774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 51078 606 51774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 52878 86090 53574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 52878 606 53574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 54678 86090 55374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 54678 606 55374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 56478 86090 57174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 56478 606 57174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 58278 86090 58974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 58278 606 58974 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 60078 86090 60774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 60078 606 60774 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 61878 86090 62574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 61878 606 62574 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 63678 86090 64374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 63678 606 64374 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 85766 65478 86090 66174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 65478 606 66174 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 282 67568 86090 67894 6 VSS
port 29 nsew ground bidirectional
rlabel metal1 s 282 282 86090 1000 6 VSS
port 29 nsew ground bidirectional
rlabel metal1 s 85372 1000 86090 67176 6 VSS
port 29 nsew ground bidirectional
rlabel metal1 s 282 1000 1000 67176 6 VSS
port 29 nsew ground bidirectional
rlabel metal1 s 282 67176 86090 67894 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 1954 26435 26070 28434 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 2249 10174 24250 11491 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27442 34494 27782 35062 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30402 65726 54622 65928 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 63926 54622 64128 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 62126 54622 62328 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 60326 54622 60528 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 58526 54622 58728 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 56726 54622 56928 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 54926 54622 55128 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 53126 54622 53328 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 51326 54622 51528 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60559 34536 60647 35387 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 58785 26435 84717 28434 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60736 10173 84482 11491 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60736 6980 84787 7595 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 82695 0 82919 1000 6 WEN[7]
port 30 nsew signal input
rlabel metal2 s 72630 0 72854 1000 6 WEN[6]
port 31 nsew signal input
rlabel metal2 s 72180 0 72404 1000 6 WEN[5]
port 32 nsew signal input
rlabel metal2 s 62115 0 62339 1000 6 WEN[4]
port 33 nsew signal input
rlabel metal2 s 23404 0 23628 1000 6 WEN[3]
port 34 nsew signal input
rlabel metal2 s 13054 0 13278 1000 6 WEN[2]
port 35 nsew signal input
rlabel metal2 s 12604 0 12828 1000 6 WEN[1]
port 36 nsew signal input
rlabel metal2 s 2539 0 2763 1000 6 WEN[0]
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 86372 68176
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2452518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2396452
<< end >>
