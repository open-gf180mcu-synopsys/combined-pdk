magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< psubdiff >>
rect 70 53483 85816 53502
rect 70 53437 89 53483
rect 135 53437 213 53483
rect 259 53437 337 53483
rect 383 53437 461 53483
rect 507 53437 585 53483
rect 631 53437 709 53483
rect 755 53437 833 53483
rect 879 53437 957 53483
rect 1003 53437 1081 53483
rect 1127 53437 1205 53483
rect 1251 53437 1329 53483
rect 1375 53437 1453 53483
rect 1499 53437 1577 53483
rect 1623 53437 1701 53483
rect 1747 53437 1825 53483
rect 1871 53437 1949 53483
rect 1995 53437 2073 53483
rect 2119 53437 2197 53483
rect 2243 53437 2321 53483
rect 2367 53437 2445 53483
rect 2491 53437 2569 53483
rect 2615 53437 2693 53483
rect 2739 53437 2817 53483
rect 2863 53437 2941 53483
rect 2987 53437 3065 53483
rect 3111 53437 3189 53483
rect 3235 53437 3313 53483
rect 3359 53437 3437 53483
rect 3483 53437 3561 53483
rect 3607 53437 3685 53483
rect 3731 53437 3809 53483
rect 3855 53437 3933 53483
rect 3979 53437 4057 53483
rect 4103 53437 4181 53483
rect 4227 53437 4305 53483
rect 4351 53437 4429 53483
rect 4475 53437 4553 53483
rect 4599 53437 4677 53483
rect 4723 53437 4801 53483
rect 4847 53437 4925 53483
rect 4971 53437 5049 53483
rect 5095 53437 5173 53483
rect 5219 53437 5297 53483
rect 5343 53437 5421 53483
rect 5467 53437 5545 53483
rect 5591 53437 5669 53483
rect 5715 53437 5793 53483
rect 5839 53437 5917 53483
rect 5963 53437 6041 53483
rect 6087 53437 6165 53483
rect 6211 53437 6289 53483
rect 6335 53437 6413 53483
rect 6459 53437 6537 53483
rect 6583 53437 6661 53483
rect 6707 53437 6785 53483
rect 6831 53437 6909 53483
rect 6955 53437 7033 53483
rect 7079 53437 7157 53483
rect 7203 53437 7281 53483
rect 7327 53437 7405 53483
rect 7451 53437 7529 53483
rect 7575 53437 7653 53483
rect 7699 53437 7777 53483
rect 7823 53437 7901 53483
rect 7947 53437 8025 53483
rect 8071 53437 8149 53483
rect 8195 53437 8273 53483
rect 8319 53437 8397 53483
rect 8443 53437 8521 53483
rect 8567 53437 8645 53483
rect 8691 53437 8769 53483
rect 8815 53437 8893 53483
rect 8939 53437 9017 53483
rect 9063 53437 9141 53483
rect 9187 53437 9265 53483
rect 9311 53437 9389 53483
rect 9435 53437 9513 53483
rect 9559 53437 9637 53483
rect 9683 53437 9761 53483
rect 9807 53437 9885 53483
rect 9931 53437 10009 53483
rect 10055 53437 10133 53483
rect 10179 53437 10257 53483
rect 10303 53437 10381 53483
rect 10427 53437 10505 53483
rect 10551 53437 10629 53483
rect 10675 53437 10753 53483
rect 10799 53437 10877 53483
rect 10923 53437 11001 53483
rect 11047 53437 11125 53483
rect 11171 53437 11249 53483
rect 11295 53437 11373 53483
rect 11419 53437 11497 53483
rect 11543 53437 11621 53483
rect 11667 53437 11745 53483
rect 11791 53437 11869 53483
rect 11915 53437 11993 53483
rect 12039 53437 12117 53483
rect 12163 53437 12241 53483
rect 12287 53437 12365 53483
rect 12411 53437 12489 53483
rect 12535 53437 12613 53483
rect 12659 53437 12737 53483
rect 12783 53437 12861 53483
rect 12907 53437 12985 53483
rect 13031 53437 13109 53483
rect 13155 53437 13233 53483
rect 13279 53437 13357 53483
rect 13403 53437 13481 53483
rect 13527 53437 13605 53483
rect 13651 53437 13729 53483
rect 13775 53437 13853 53483
rect 13899 53437 13977 53483
rect 14023 53437 14101 53483
rect 14147 53437 14225 53483
rect 14271 53437 14349 53483
rect 14395 53437 14473 53483
rect 14519 53437 14597 53483
rect 14643 53437 14721 53483
rect 14767 53437 14845 53483
rect 14891 53437 14969 53483
rect 15015 53437 15093 53483
rect 15139 53437 15217 53483
rect 15263 53437 15341 53483
rect 15387 53437 15465 53483
rect 15511 53437 15589 53483
rect 15635 53437 15713 53483
rect 15759 53437 15837 53483
rect 15883 53437 15961 53483
rect 16007 53437 16085 53483
rect 16131 53437 16209 53483
rect 16255 53437 16333 53483
rect 16379 53437 16457 53483
rect 16503 53437 16581 53483
rect 16627 53437 16705 53483
rect 16751 53437 16829 53483
rect 16875 53437 16953 53483
rect 16999 53437 17077 53483
rect 17123 53437 17201 53483
rect 17247 53437 17325 53483
rect 17371 53437 17449 53483
rect 17495 53437 17573 53483
rect 17619 53437 17697 53483
rect 17743 53437 17821 53483
rect 17867 53437 17945 53483
rect 17991 53437 18069 53483
rect 18115 53437 18193 53483
rect 18239 53437 18317 53483
rect 18363 53437 18441 53483
rect 18487 53437 18565 53483
rect 18611 53437 18689 53483
rect 18735 53437 18813 53483
rect 18859 53437 18937 53483
rect 18983 53437 19061 53483
rect 19107 53437 19185 53483
rect 19231 53437 19309 53483
rect 19355 53437 19433 53483
rect 19479 53437 19557 53483
rect 19603 53437 19681 53483
rect 19727 53437 19805 53483
rect 19851 53437 19929 53483
rect 19975 53437 20053 53483
rect 20099 53437 20177 53483
rect 20223 53437 20301 53483
rect 20347 53437 20425 53483
rect 20471 53437 20549 53483
rect 20595 53437 20673 53483
rect 20719 53437 20797 53483
rect 20843 53437 20921 53483
rect 20967 53437 21045 53483
rect 21091 53437 21169 53483
rect 21215 53437 21293 53483
rect 21339 53437 21417 53483
rect 21463 53437 21541 53483
rect 21587 53437 21665 53483
rect 21711 53437 21789 53483
rect 21835 53437 21913 53483
rect 21959 53437 22037 53483
rect 22083 53437 22161 53483
rect 22207 53437 22285 53483
rect 22331 53437 22409 53483
rect 22455 53437 22533 53483
rect 22579 53437 22657 53483
rect 22703 53437 22781 53483
rect 22827 53437 22905 53483
rect 22951 53437 23029 53483
rect 23075 53437 23153 53483
rect 23199 53437 23277 53483
rect 23323 53437 23401 53483
rect 23447 53437 23525 53483
rect 23571 53437 23649 53483
rect 23695 53437 23773 53483
rect 23819 53437 23897 53483
rect 23943 53437 24021 53483
rect 24067 53437 24145 53483
rect 24191 53437 24269 53483
rect 24315 53437 24393 53483
rect 24439 53437 24517 53483
rect 24563 53437 24641 53483
rect 24687 53437 24765 53483
rect 24811 53437 24889 53483
rect 24935 53437 25013 53483
rect 25059 53437 25137 53483
rect 25183 53437 25261 53483
rect 25307 53437 25385 53483
rect 25431 53437 25509 53483
rect 25555 53437 25633 53483
rect 25679 53437 25757 53483
rect 25803 53437 25881 53483
rect 25927 53437 26005 53483
rect 26051 53437 26129 53483
rect 26175 53437 26253 53483
rect 26299 53437 26377 53483
rect 26423 53437 26501 53483
rect 26547 53437 26625 53483
rect 26671 53437 26749 53483
rect 26795 53437 26873 53483
rect 26919 53437 26997 53483
rect 27043 53437 27121 53483
rect 27167 53437 27245 53483
rect 27291 53437 27369 53483
rect 27415 53437 27493 53483
rect 27539 53437 27617 53483
rect 27663 53437 27741 53483
rect 27787 53437 27865 53483
rect 27911 53437 27989 53483
rect 28035 53437 28113 53483
rect 28159 53437 28237 53483
rect 28283 53437 28361 53483
rect 28407 53437 28485 53483
rect 28531 53437 28609 53483
rect 28655 53437 28733 53483
rect 28779 53437 28857 53483
rect 28903 53437 28981 53483
rect 29027 53437 29105 53483
rect 29151 53437 29229 53483
rect 29275 53437 29353 53483
rect 29399 53437 29477 53483
rect 29523 53437 29601 53483
rect 29647 53437 29725 53483
rect 29771 53437 29849 53483
rect 29895 53437 29973 53483
rect 30019 53437 30097 53483
rect 30143 53437 30221 53483
rect 30267 53437 30345 53483
rect 30391 53437 30469 53483
rect 30515 53437 30593 53483
rect 30639 53437 30717 53483
rect 30763 53437 30841 53483
rect 30887 53437 30965 53483
rect 31011 53437 31089 53483
rect 31135 53437 31213 53483
rect 31259 53437 31337 53483
rect 31383 53437 31461 53483
rect 31507 53437 31585 53483
rect 31631 53437 31709 53483
rect 31755 53437 31833 53483
rect 31879 53437 31957 53483
rect 32003 53437 32081 53483
rect 32127 53437 32205 53483
rect 32251 53437 32329 53483
rect 32375 53437 32453 53483
rect 32499 53437 32577 53483
rect 32623 53437 32701 53483
rect 32747 53437 32825 53483
rect 32871 53437 32949 53483
rect 32995 53437 33073 53483
rect 33119 53437 33197 53483
rect 33243 53437 33321 53483
rect 33367 53437 33445 53483
rect 33491 53437 33569 53483
rect 33615 53437 33693 53483
rect 33739 53437 33817 53483
rect 33863 53437 33941 53483
rect 33987 53437 34065 53483
rect 34111 53437 34189 53483
rect 34235 53437 34313 53483
rect 34359 53437 34437 53483
rect 34483 53437 34561 53483
rect 34607 53437 34685 53483
rect 34731 53437 34809 53483
rect 34855 53437 34933 53483
rect 34979 53437 35057 53483
rect 35103 53437 35181 53483
rect 35227 53437 35305 53483
rect 35351 53437 35429 53483
rect 35475 53437 35553 53483
rect 35599 53437 35677 53483
rect 35723 53437 35801 53483
rect 35847 53437 35925 53483
rect 35971 53437 36049 53483
rect 36095 53437 36173 53483
rect 36219 53437 36297 53483
rect 36343 53437 36421 53483
rect 36467 53437 36545 53483
rect 36591 53437 36669 53483
rect 36715 53437 36793 53483
rect 36839 53437 36917 53483
rect 36963 53437 37041 53483
rect 37087 53437 37165 53483
rect 37211 53437 37289 53483
rect 37335 53437 37413 53483
rect 37459 53437 37537 53483
rect 37583 53437 37661 53483
rect 37707 53437 37785 53483
rect 37831 53437 37909 53483
rect 37955 53437 38033 53483
rect 38079 53437 38157 53483
rect 38203 53437 38281 53483
rect 38327 53437 38405 53483
rect 38451 53437 38529 53483
rect 38575 53437 38653 53483
rect 38699 53437 38777 53483
rect 38823 53437 38901 53483
rect 38947 53437 39025 53483
rect 39071 53437 39149 53483
rect 39195 53437 39273 53483
rect 39319 53437 39397 53483
rect 39443 53437 39521 53483
rect 39567 53437 39645 53483
rect 39691 53437 39769 53483
rect 39815 53437 39893 53483
rect 39939 53437 40017 53483
rect 40063 53437 40141 53483
rect 40187 53437 40265 53483
rect 40311 53437 40389 53483
rect 40435 53437 40513 53483
rect 40559 53437 40637 53483
rect 40683 53437 40761 53483
rect 40807 53437 40885 53483
rect 40931 53437 41009 53483
rect 41055 53437 41133 53483
rect 41179 53437 41257 53483
rect 41303 53437 41381 53483
rect 41427 53437 41505 53483
rect 41551 53437 41629 53483
rect 41675 53437 41753 53483
rect 41799 53437 41877 53483
rect 41923 53437 42001 53483
rect 42047 53437 42125 53483
rect 42171 53437 42249 53483
rect 42295 53437 42373 53483
rect 42419 53437 42497 53483
rect 42543 53437 42621 53483
rect 42667 53437 42745 53483
rect 42791 53437 42869 53483
rect 42915 53437 42993 53483
rect 43039 53437 43117 53483
rect 43163 53437 43241 53483
rect 43287 53437 43365 53483
rect 43411 53437 43489 53483
rect 43535 53437 43613 53483
rect 43659 53437 43737 53483
rect 43783 53437 43861 53483
rect 43907 53437 43985 53483
rect 44031 53437 44109 53483
rect 44155 53437 44233 53483
rect 44279 53437 44357 53483
rect 44403 53437 44481 53483
rect 44527 53437 44605 53483
rect 44651 53437 44729 53483
rect 44775 53437 44853 53483
rect 44899 53437 44977 53483
rect 45023 53437 45101 53483
rect 45147 53437 45225 53483
rect 45271 53437 45349 53483
rect 45395 53437 45473 53483
rect 45519 53437 45597 53483
rect 45643 53437 45721 53483
rect 45767 53437 45845 53483
rect 45891 53437 45969 53483
rect 46015 53437 46093 53483
rect 46139 53437 46217 53483
rect 46263 53437 46341 53483
rect 46387 53437 46465 53483
rect 46511 53437 46589 53483
rect 46635 53437 46713 53483
rect 46759 53437 46837 53483
rect 46883 53437 46961 53483
rect 47007 53437 47085 53483
rect 47131 53437 47209 53483
rect 47255 53437 47333 53483
rect 47379 53437 47457 53483
rect 47503 53437 47581 53483
rect 47627 53437 47705 53483
rect 47751 53437 47829 53483
rect 47875 53437 47953 53483
rect 47999 53437 48077 53483
rect 48123 53437 48201 53483
rect 48247 53437 48325 53483
rect 48371 53437 48449 53483
rect 48495 53437 48573 53483
rect 48619 53437 48697 53483
rect 48743 53437 48821 53483
rect 48867 53437 48945 53483
rect 48991 53437 49069 53483
rect 49115 53437 49193 53483
rect 49239 53437 49317 53483
rect 49363 53437 49441 53483
rect 49487 53437 49565 53483
rect 49611 53437 49689 53483
rect 49735 53437 49813 53483
rect 49859 53437 49937 53483
rect 49983 53437 50061 53483
rect 50107 53437 50185 53483
rect 50231 53437 50309 53483
rect 50355 53437 50433 53483
rect 50479 53437 50557 53483
rect 50603 53437 50681 53483
rect 50727 53437 50805 53483
rect 50851 53437 50929 53483
rect 50975 53437 51053 53483
rect 51099 53437 51177 53483
rect 51223 53437 51301 53483
rect 51347 53437 51425 53483
rect 51471 53437 51549 53483
rect 51595 53437 51673 53483
rect 51719 53437 51797 53483
rect 51843 53437 51921 53483
rect 51967 53437 52045 53483
rect 52091 53437 52169 53483
rect 52215 53437 52293 53483
rect 52339 53437 52417 53483
rect 52463 53437 52541 53483
rect 52587 53437 52665 53483
rect 52711 53437 52789 53483
rect 52835 53437 52913 53483
rect 52959 53437 53037 53483
rect 53083 53437 53161 53483
rect 53207 53437 53285 53483
rect 53331 53437 53409 53483
rect 53455 53437 53533 53483
rect 53579 53437 53657 53483
rect 53703 53437 53781 53483
rect 53827 53437 53905 53483
rect 53951 53437 54029 53483
rect 54075 53437 54153 53483
rect 54199 53437 54277 53483
rect 54323 53437 54401 53483
rect 54447 53437 54525 53483
rect 54571 53437 54649 53483
rect 54695 53437 54773 53483
rect 54819 53437 54897 53483
rect 54943 53437 55021 53483
rect 55067 53437 55145 53483
rect 55191 53437 55269 53483
rect 55315 53437 55393 53483
rect 55439 53437 55517 53483
rect 55563 53437 55641 53483
rect 55687 53437 55765 53483
rect 55811 53437 55889 53483
rect 55935 53437 56013 53483
rect 56059 53437 56137 53483
rect 56183 53437 56261 53483
rect 56307 53437 56385 53483
rect 56431 53437 56509 53483
rect 56555 53437 56633 53483
rect 56679 53437 56757 53483
rect 56803 53437 56881 53483
rect 56927 53437 57005 53483
rect 57051 53437 57129 53483
rect 57175 53437 57253 53483
rect 57299 53437 57377 53483
rect 57423 53437 57501 53483
rect 57547 53437 57625 53483
rect 57671 53437 57749 53483
rect 57795 53437 57873 53483
rect 57919 53437 57997 53483
rect 58043 53437 58121 53483
rect 58167 53437 58245 53483
rect 58291 53437 58369 53483
rect 58415 53437 58493 53483
rect 58539 53437 58617 53483
rect 58663 53437 58741 53483
rect 58787 53437 58865 53483
rect 58911 53437 58989 53483
rect 59035 53437 59113 53483
rect 59159 53437 59237 53483
rect 59283 53437 59361 53483
rect 59407 53437 59485 53483
rect 59531 53437 59609 53483
rect 59655 53437 59733 53483
rect 59779 53437 59857 53483
rect 59903 53437 59981 53483
rect 60027 53437 60105 53483
rect 60151 53437 60229 53483
rect 60275 53437 60353 53483
rect 60399 53437 60477 53483
rect 60523 53437 60601 53483
rect 60647 53437 60725 53483
rect 60771 53437 60849 53483
rect 60895 53437 60973 53483
rect 61019 53437 61097 53483
rect 61143 53437 61221 53483
rect 61267 53437 61345 53483
rect 61391 53437 61469 53483
rect 61515 53437 61593 53483
rect 61639 53437 61717 53483
rect 61763 53437 61841 53483
rect 61887 53437 61965 53483
rect 62011 53437 62089 53483
rect 62135 53437 62213 53483
rect 62259 53437 62337 53483
rect 62383 53437 62461 53483
rect 62507 53437 62585 53483
rect 62631 53437 62709 53483
rect 62755 53437 62833 53483
rect 62879 53437 62957 53483
rect 63003 53437 63081 53483
rect 63127 53437 63205 53483
rect 63251 53437 63329 53483
rect 63375 53437 63453 53483
rect 63499 53437 63577 53483
rect 63623 53437 63701 53483
rect 63747 53437 63825 53483
rect 63871 53437 63949 53483
rect 63995 53437 64073 53483
rect 64119 53437 64197 53483
rect 64243 53437 64321 53483
rect 64367 53437 64445 53483
rect 64491 53437 64569 53483
rect 64615 53437 64693 53483
rect 64739 53437 64817 53483
rect 64863 53437 64941 53483
rect 64987 53437 65065 53483
rect 65111 53437 65189 53483
rect 65235 53437 65313 53483
rect 65359 53437 65437 53483
rect 65483 53437 65561 53483
rect 65607 53437 65685 53483
rect 65731 53437 65809 53483
rect 65855 53437 65933 53483
rect 65979 53437 66057 53483
rect 66103 53437 66181 53483
rect 66227 53437 66305 53483
rect 66351 53437 66429 53483
rect 66475 53437 66553 53483
rect 66599 53437 66677 53483
rect 66723 53437 66801 53483
rect 66847 53437 66925 53483
rect 66971 53437 67049 53483
rect 67095 53437 67173 53483
rect 67219 53437 67297 53483
rect 67343 53437 67421 53483
rect 67467 53437 67545 53483
rect 67591 53437 67669 53483
rect 67715 53437 67793 53483
rect 67839 53437 67917 53483
rect 67963 53437 68041 53483
rect 68087 53437 68165 53483
rect 68211 53437 68289 53483
rect 68335 53437 68413 53483
rect 68459 53437 68537 53483
rect 68583 53437 68661 53483
rect 68707 53437 68785 53483
rect 68831 53437 68909 53483
rect 68955 53437 69033 53483
rect 69079 53437 69157 53483
rect 69203 53437 69281 53483
rect 69327 53437 69405 53483
rect 69451 53437 69529 53483
rect 69575 53437 69653 53483
rect 69699 53437 69777 53483
rect 69823 53437 69901 53483
rect 69947 53437 70025 53483
rect 70071 53437 70149 53483
rect 70195 53437 70273 53483
rect 70319 53437 70397 53483
rect 70443 53437 70521 53483
rect 70567 53437 70645 53483
rect 70691 53437 70769 53483
rect 70815 53437 70893 53483
rect 70939 53437 71017 53483
rect 71063 53437 71141 53483
rect 71187 53437 71265 53483
rect 71311 53437 71389 53483
rect 71435 53437 71513 53483
rect 71559 53437 71637 53483
rect 71683 53437 71761 53483
rect 71807 53437 71885 53483
rect 71931 53437 72009 53483
rect 72055 53437 72133 53483
rect 72179 53437 72257 53483
rect 72303 53437 72381 53483
rect 72427 53437 72505 53483
rect 72551 53437 72629 53483
rect 72675 53437 72753 53483
rect 72799 53437 72877 53483
rect 72923 53437 73001 53483
rect 73047 53437 73125 53483
rect 73171 53437 73249 53483
rect 73295 53437 73373 53483
rect 73419 53437 73497 53483
rect 73543 53437 73621 53483
rect 73667 53437 73745 53483
rect 73791 53437 73869 53483
rect 73915 53437 73993 53483
rect 74039 53437 74117 53483
rect 74163 53437 74241 53483
rect 74287 53437 74365 53483
rect 74411 53437 74489 53483
rect 74535 53437 74613 53483
rect 74659 53437 74737 53483
rect 74783 53437 74861 53483
rect 74907 53437 74985 53483
rect 75031 53437 75109 53483
rect 75155 53437 75233 53483
rect 75279 53437 75357 53483
rect 75403 53437 75481 53483
rect 75527 53437 75605 53483
rect 75651 53437 75729 53483
rect 75775 53437 75853 53483
rect 75899 53437 75977 53483
rect 76023 53437 76101 53483
rect 76147 53437 76225 53483
rect 76271 53437 76349 53483
rect 76395 53437 76473 53483
rect 76519 53437 76597 53483
rect 76643 53437 76721 53483
rect 76767 53437 76845 53483
rect 76891 53437 76969 53483
rect 77015 53437 77093 53483
rect 77139 53437 77217 53483
rect 77263 53437 77341 53483
rect 77387 53437 77465 53483
rect 77511 53437 77589 53483
rect 77635 53437 77713 53483
rect 77759 53437 77837 53483
rect 77883 53437 77961 53483
rect 78007 53437 78085 53483
rect 78131 53437 78209 53483
rect 78255 53437 78333 53483
rect 78379 53437 78457 53483
rect 78503 53437 78581 53483
rect 78627 53437 78705 53483
rect 78751 53437 78829 53483
rect 78875 53437 78953 53483
rect 78999 53437 79077 53483
rect 79123 53437 79201 53483
rect 79247 53437 79325 53483
rect 79371 53437 79449 53483
rect 79495 53437 79573 53483
rect 79619 53437 79697 53483
rect 79743 53437 79821 53483
rect 79867 53437 79945 53483
rect 79991 53437 80069 53483
rect 80115 53437 80193 53483
rect 80239 53437 80317 53483
rect 80363 53437 80441 53483
rect 80487 53437 80565 53483
rect 80611 53437 80689 53483
rect 80735 53437 80813 53483
rect 80859 53437 80937 53483
rect 80983 53437 81061 53483
rect 81107 53437 81185 53483
rect 81231 53437 81309 53483
rect 81355 53437 81433 53483
rect 81479 53437 81557 53483
rect 81603 53437 81681 53483
rect 81727 53437 81805 53483
rect 81851 53437 81929 53483
rect 81975 53437 82053 53483
rect 82099 53437 82177 53483
rect 82223 53437 82301 53483
rect 82347 53437 82425 53483
rect 82471 53437 82549 53483
rect 82595 53437 82673 53483
rect 82719 53437 82797 53483
rect 82843 53437 82921 53483
rect 82967 53437 83045 53483
rect 83091 53437 83169 53483
rect 83215 53437 83293 53483
rect 83339 53437 83417 53483
rect 83463 53437 83541 53483
rect 83587 53437 83665 53483
rect 83711 53437 83789 53483
rect 83835 53437 83913 53483
rect 83959 53437 84037 53483
rect 84083 53437 84161 53483
rect 84207 53437 84285 53483
rect 84331 53437 84409 53483
rect 84455 53437 84533 53483
rect 84579 53437 84657 53483
rect 84703 53437 84781 53483
rect 84827 53437 84905 53483
rect 84951 53437 85029 53483
rect 85075 53437 85153 53483
rect 85199 53437 85277 53483
rect 85323 53437 85401 53483
rect 85447 53437 85525 53483
rect 85571 53437 85649 53483
rect 85695 53437 85816 53483
rect 70 53359 85816 53437
rect 70 53313 89 53359
rect 135 53313 213 53359
rect 259 53313 337 53359
rect 383 53313 461 53359
rect 507 53313 585 53359
rect 631 53313 709 53359
rect 755 53313 833 53359
rect 879 53313 957 53359
rect 1003 53313 1081 53359
rect 1127 53313 1205 53359
rect 1251 53313 1329 53359
rect 1375 53313 1453 53359
rect 1499 53313 1577 53359
rect 1623 53313 1701 53359
rect 1747 53313 1825 53359
rect 1871 53313 1949 53359
rect 1995 53313 2073 53359
rect 2119 53313 2197 53359
rect 2243 53313 2321 53359
rect 2367 53313 2445 53359
rect 2491 53313 2569 53359
rect 2615 53313 2693 53359
rect 2739 53313 2817 53359
rect 2863 53313 2941 53359
rect 2987 53313 3065 53359
rect 3111 53313 3189 53359
rect 3235 53313 3313 53359
rect 3359 53313 3437 53359
rect 3483 53313 3561 53359
rect 3607 53313 3685 53359
rect 3731 53313 3809 53359
rect 3855 53313 3933 53359
rect 3979 53313 4057 53359
rect 4103 53313 4181 53359
rect 4227 53313 4305 53359
rect 4351 53313 4429 53359
rect 4475 53313 4553 53359
rect 4599 53313 4677 53359
rect 4723 53313 4801 53359
rect 4847 53313 4925 53359
rect 4971 53313 5049 53359
rect 5095 53313 5173 53359
rect 5219 53313 5297 53359
rect 5343 53313 5421 53359
rect 5467 53313 5545 53359
rect 5591 53313 5669 53359
rect 5715 53313 5793 53359
rect 5839 53313 5917 53359
rect 5963 53313 6041 53359
rect 6087 53313 6165 53359
rect 6211 53313 6289 53359
rect 6335 53313 6413 53359
rect 6459 53313 6537 53359
rect 6583 53313 6661 53359
rect 6707 53313 6785 53359
rect 6831 53313 6909 53359
rect 6955 53313 7033 53359
rect 7079 53313 7157 53359
rect 7203 53313 7281 53359
rect 7327 53313 7405 53359
rect 7451 53313 7529 53359
rect 7575 53313 7653 53359
rect 7699 53313 7777 53359
rect 7823 53313 7901 53359
rect 7947 53313 8025 53359
rect 8071 53313 8149 53359
rect 8195 53313 8273 53359
rect 8319 53313 8397 53359
rect 8443 53313 8521 53359
rect 8567 53313 8645 53359
rect 8691 53313 8769 53359
rect 8815 53313 8893 53359
rect 8939 53313 9017 53359
rect 9063 53313 9141 53359
rect 9187 53313 9265 53359
rect 9311 53313 9389 53359
rect 9435 53313 9513 53359
rect 9559 53313 9637 53359
rect 9683 53313 9761 53359
rect 9807 53313 9885 53359
rect 9931 53313 10009 53359
rect 10055 53313 10133 53359
rect 10179 53313 10257 53359
rect 10303 53313 10381 53359
rect 10427 53313 10505 53359
rect 10551 53313 10629 53359
rect 10675 53313 10753 53359
rect 10799 53313 10877 53359
rect 10923 53313 11001 53359
rect 11047 53313 11125 53359
rect 11171 53313 11249 53359
rect 11295 53313 11373 53359
rect 11419 53313 11497 53359
rect 11543 53313 11621 53359
rect 11667 53313 11745 53359
rect 11791 53313 11869 53359
rect 11915 53313 11993 53359
rect 12039 53313 12117 53359
rect 12163 53313 12241 53359
rect 12287 53313 12365 53359
rect 12411 53313 12489 53359
rect 12535 53313 12613 53359
rect 12659 53313 12737 53359
rect 12783 53313 12861 53359
rect 12907 53313 12985 53359
rect 13031 53313 13109 53359
rect 13155 53313 13233 53359
rect 13279 53313 13357 53359
rect 13403 53313 13481 53359
rect 13527 53313 13605 53359
rect 13651 53313 13729 53359
rect 13775 53313 13853 53359
rect 13899 53313 13977 53359
rect 14023 53313 14101 53359
rect 14147 53313 14225 53359
rect 14271 53313 14349 53359
rect 14395 53313 14473 53359
rect 14519 53313 14597 53359
rect 14643 53313 14721 53359
rect 14767 53313 14845 53359
rect 14891 53313 14969 53359
rect 15015 53313 15093 53359
rect 15139 53313 15217 53359
rect 15263 53313 15341 53359
rect 15387 53313 15465 53359
rect 15511 53313 15589 53359
rect 15635 53313 15713 53359
rect 15759 53313 15837 53359
rect 15883 53313 15961 53359
rect 16007 53313 16085 53359
rect 16131 53313 16209 53359
rect 16255 53313 16333 53359
rect 16379 53313 16457 53359
rect 16503 53313 16581 53359
rect 16627 53313 16705 53359
rect 16751 53313 16829 53359
rect 16875 53313 16953 53359
rect 16999 53313 17077 53359
rect 17123 53313 17201 53359
rect 17247 53313 17325 53359
rect 17371 53313 17449 53359
rect 17495 53313 17573 53359
rect 17619 53313 17697 53359
rect 17743 53313 17821 53359
rect 17867 53313 17945 53359
rect 17991 53313 18069 53359
rect 18115 53313 18193 53359
rect 18239 53313 18317 53359
rect 18363 53313 18441 53359
rect 18487 53313 18565 53359
rect 18611 53313 18689 53359
rect 18735 53313 18813 53359
rect 18859 53313 18937 53359
rect 18983 53313 19061 53359
rect 19107 53313 19185 53359
rect 19231 53313 19309 53359
rect 19355 53313 19433 53359
rect 19479 53313 19557 53359
rect 19603 53313 19681 53359
rect 19727 53313 19805 53359
rect 19851 53313 19929 53359
rect 19975 53313 20053 53359
rect 20099 53313 20177 53359
rect 20223 53313 20301 53359
rect 20347 53313 20425 53359
rect 20471 53313 20549 53359
rect 20595 53313 20673 53359
rect 20719 53313 20797 53359
rect 20843 53313 20921 53359
rect 20967 53313 21045 53359
rect 21091 53313 21169 53359
rect 21215 53313 21293 53359
rect 21339 53313 21417 53359
rect 21463 53313 21541 53359
rect 21587 53313 21665 53359
rect 21711 53313 21789 53359
rect 21835 53313 21913 53359
rect 21959 53313 22037 53359
rect 22083 53313 22161 53359
rect 22207 53313 22285 53359
rect 22331 53313 22409 53359
rect 22455 53313 22533 53359
rect 22579 53313 22657 53359
rect 22703 53313 22781 53359
rect 22827 53313 22905 53359
rect 22951 53313 23029 53359
rect 23075 53313 23153 53359
rect 23199 53313 23277 53359
rect 23323 53313 23401 53359
rect 23447 53313 23525 53359
rect 23571 53313 23649 53359
rect 23695 53313 23773 53359
rect 23819 53313 23897 53359
rect 23943 53313 24021 53359
rect 24067 53313 24145 53359
rect 24191 53313 24269 53359
rect 24315 53313 24393 53359
rect 24439 53313 24517 53359
rect 24563 53313 24641 53359
rect 24687 53313 24765 53359
rect 24811 53313 24889 53359
rect 24935 53313 25013 53359
rect 25059 53313 25137 53359
rect 25183 53313 25261 53359
rect 25307 53313 25385 53359
rect 25431 53313 25509 53359
rect 25555 53313 25633 53359
rect 25679 53313 25757 53359
rect 25803 53313 25881 53359
rect 25927 53313 26005 53359
rect 26051 53313 26129 53359
rect 26175 53313 26253 53359
rect 26299 53313 26377 53359
rect 26423 53313 26501 53359
rect 26547 53313 26625 53359
rect 26671 53313 26749 53359
rect 26795 53313 26873 53359
rect 26919 53313 26997 53359
rect 27043 53313 27121 53359
rect 27167 53313 27245 53359
rect 27291 53313 27369 53359
rect 27415 53313 27493 53359
rect 27539 53313 27617 53359
rect 27663 53313 27741 53359
rect 27787 53313 27865 53359
rect 27911 53313 27989 53359
rect 28035 53313 28113 53359
rect 28159 53313 28237 53359
rect 28283 53313 28361 53359
rect 28407 53313 28485 53359
rect 28531 53313 28609 53359
rect 28655 53313 28733 53359
rect 28779 53313 28857 53359
rect 28903 53313 28981 53359
rect 29027 53313 29105 53359
rect 29151 53313 29229 53359
rect 29275 53313 29353 53359
rect 29399 53313 29477 53359
rect 29523 53313 29601 53359
rect 29647 53313 29725 53359
rect 29771 53313 29849 53359
rect 29895 53313 29973 53359
rect 30019 53313 30097 53359
rect 30143 53313 30221 53359
rect 30267 53313 30345 53359
rect 30391 53313 30469 53359
rect 30515 53313 30593 53359
rect 30639 53313 30717 53359
rect 30763 53313 30841 53359
rect 30887 53313 30965 53359
rect 31011 53313 31089 53359
rect 31135 53313 31213 53359
rect 31259 53313 31337 53359
rect 31383 53313 31461 53359
rect 31507 53313 31585 53359
rect 31631 53313 31709 53359
rect 31755 53313 31833 53359
rect 31879 53313 31957 53359
rect 32003 53313 32081 53359
rect 32127 53313 32205 53359
rect 32251 53313 32329 53359
rect 32375 53313 32453 53359
rect 32499 53313 32577 53359
rect 32623 53313 32701 53359
rect 32747 53313 32825 53359
rect 32871 53313 32949 53359
rect 32995 53313 33073 53359
rect 33119 53313 33197 53359
rect 33243 53313 33321 53359
rect 33367 53313 33445 53359
rect 33491 53313 33569 53359
rect 33615 53313 33693 53359
rect 33739 53313 33817 53359
rect 33863 53313 33941 53359
rect 33987 53313 34065 53359
rect 34111 53313 34189 53359
rect 34235 53313 34313 53359
rect 34359 53313 34437 53359
rect 34483 53313 34561 53359
rect 34607 53313 34685 53359
rect 34731 53313 34809 53359
rect 34855 53313 34933 53359
rect 34979 53313 35057 53359
rect 35103 53313 35181 53359
rect 35227 53313 35305 53359
rect 35351 53313 35429 53359
rect 35475 53313 35553 53359
rect 35599 53313 35677 53359
rect 35723 53313 35801 53359
rect 35847 53313 35925 53359
rect 35971 53313 36049 53359
rect 36095 53313 36173 53359
rect 36219 53313 36297 53359
rect 36343 53313 36421 53359
rect 36467 53313 36545 53359
rect 36591 53313 36669 53359
rect 36715 53313 36793 53359
rect 36839 53313 36917 53359
rect 36963 53313 37041 53359
rect 37087 53313 37165 53359
rect 37211 53313 37289 53359
rect 37335 53313 37413 53359
rect 37459 53313 37537 53359
rect 37583 53313 37661 53359
rect 37707 53313 37785 53359
rect 37831 53313 37909 53359
rect 37955 53313 38033 53359
rect 38079 53313 38157 53359
rect 38203 53313 38281 53359
rect 38327 53313 38405 53359
rect 38451 53313 38529 53359
rect 38575 53313 38653 53359
rect 38699 53313 38777 53359
rect 38823 53313 38901 53359
rect 38947 53313 39025 53359
rect 39071 53313 39149 53359
rect 39195 53313 39273 53359
rect 39319 53313 39397 53359
rect 39443 53313 39521 53359
rect 39567 53313 39645 53359
rect 39691 53313 39769 53359
rect 39815 53313 39893 53359
rect 39939 53313 40017 53359
rect 40063 53313 40141 53359
rect 40187 53313 40265 53359
rect 40311 53313 40389 53359
rect 40435 53313 40513 53359
rect 40559 53313 40637 53359
rect 40683 53313 40761 53359
rect 40807 53313 40885 53359
rect 40931 53313 41009 53359
rect 41055 53313 41133 53359
rect 41179 53313 41257 53359
rect 41303 53313 41381 53359
rect 41427 53313 41505 53359
rect 41551 53313 41629 53359
rect 41675 53313 41753 53359
rect 41799 53313 41877 53359
rect 41923 53313 42001 53359
rect 42047 53313 42125 53359
rect 42171 53313 42249 53359
rect 42295 53313 42373 53359
rect 42419 53313 42497 53359
rect 42543 53313 42621 53359
rect 42667 53313 42745 53359
rect 42791 53313 42869 53359
rect 42915 53313 42993 53359
rect 43039 53313 43117 53359
rect 43163 53313 43241 53359
rect 43287 53313 43365 53359
rect 43411 53313 43489 53359
rect 43535 53313 43613 53359
rect 43659 53313 43737 53359
rect 43783 53313 43861 53359
rect 43907 53313 43985 53359
rect 44031 53313 44109 53359
rect 44155 53313 44233 53359
rect 44279 53313 44357 53359
rect 44403 53313 44481 53359
rect 44527 53313 44605 53359
rect 44651 53313 44729 53359
rect 44775 53313 44853 53359
rect 44899 53313 44977 53359
rect 45023 53313 45101 53359
rect 45147 53313 45225 53359
rect 45271 53313 45349 53359
rect 45395 53313 45473 53359
rect 45519 53313 45597 53359
rect 45643 53313 45721 53359
rect 45767 53313 45845 53359
rect 45891 53313 45969 53359
rect 46015 53313 46093 53359
rect 46139 53313 46217 53359
rect 46263 53313 46341 53359
rect 46387 53313 46465 53359
rect 46511 53313 46589 53359
rect 46635 53313 46713 53359
rect 46759 53313 46837 53359
rect 46883 53313 46961 53359
rect 47007 53313 47085 53359
rect 47131 53313 47209 53359
rect 47255 53313 47333 53359
rect 47379 53313 47457 53359
rect 47503 53313 47581 53359
rect 47627 53313 47705 53359
rect 47751 53313 47829 53359
rect 47875 53313 47953 53359
rect 47999 53313 48077 53359
rect 48123 53313 48201 53359
rect 48247 53313 48325 53359
rect 48371 53313 48449 53359
rect 48495 53313 48573 53359
rect 48619 53313 48697 53359
rect 48743 53313 48821 53359
rect 48867 53313 48945 53359
rect 48991 53313 49069 53359
rect 49115 53313 49193 53359
rect 49239 53313 49317 53359
rect 49363 53313 49441 53359
rect 49487 53313 49565 53359
rect 49611 53313 49689 53359
rect 49735 53313 49813 53359
rect 49859 53313 49937 53359
rect 49983 53313 50061 53359
rect 50107 53313 50185 53359
rect 50231 53313 50309 53359
rect 50355 53313 50433 53359
rect 50479 53313 50557 53359
rect 50603 53313 50681 53359
rect 50727 53313 50805 53359
rect 50851 53313 50929 53359
rect 50975 53313 51053 53359
rect 51099 53313 51177 53359
rect 51223 53313 51301 53359
rect 51347 53313 51425 53359
rect 51471 53313 51549 53359
rect 51595 53313 51673 53359
rect 51719 53313 51797 53359
rect 51843 53313 51921 53359
rect 51967 53313 52045 53359
rect 52091 53313 52169 53359
rect 52215 53313 52293 53359
rect 52339 53313 52417 53359
rect 52463 53313 52541 53359
rect 52587 53313 52665 53359
rect 52711 53313 52789 53359
rect 52835 53313 52913 53359
rect 52959 53313 53037 53359
rect 53083 53313 53161 53359
rect 53207 53313 53285 53359
rect 53331 53313 53409 53359
rect 53455 53313 53533 53359
rect 53579 53313 53657 53359
rect 53703 53313 53781 53359
rect 53827 53313 53905 53359
rect 53951 53313 54029 53359
rect 54075 53313 54153 53359
rect 54199 53313 54277 53359
rect 54323 53313 54401 53359
rect 54447 53313 54525 53359
rect 54571 53313 54649 53359
rect 54695 53313 54773 53359
rect 54819 53313 54897 53359
rect 54943 53313 55021 53359
rect 55067 53313 55145 53359
rect 55191 53313 55269 53359
rect 55315 53313 55393 53359
rect 55439 53313 55517 53359
rect 55563 53313 55641 53359
rect 55687 53313 55765 53359
rect 55811 53313 55889 53359
rect 55935 53313 56013 53359
rect 56059 53313 56137 53359
rect 56183 53313 56261 53359
rect 56307 53313 56385 53359
rect 56431 53313 56509 53359
rect 56555 53313 56633 53359
rect 56679 53313 56757 53359
rect 56803 53313 56881 53359
rect 56927 53313 57005 53359
rect 57051 53313 57129 53359
rect 57175 53313 57253 53359
rect 57299 53313 57377 53359
rect 57423 53313 57501 53359
rect 57547 53313 57625 53359
rect 57671 53313 57749 53359
rect 57795 53313 57873 53359
rect 57919 53313 57997 53359
rect 58043 53313 58121 53359
rect 58167 53313 58245 53359
rect 58291 53313 58369 53359
rect 58415 53313 58493 53359
rect 58539 53313 58617 53359
rect 58663 53313 58741 53359
rect 58787 53313 58865 53359
rect 58911 53313 58989 53359
rect 59035 53313 59113 53359
rect 59159 53313 59237 53359
rect 59283 53313 59361 53359
rect 59407 53313 59485 53359
rect 59531 53313 59609 53359
rect 59655 53313 59733 53359
rect 59779 53313 59857 53359
rect 59903 53313 59981 53359
rect 60027 53313 60105 53359
rect 60151 53313 60229 53359
rect 60275 53313 60353 53359
rect 60399 53313 60477 53359
rect 60523 53313 60601 53359
rect 60647 53313 60725 53359
rect 60771 53313 60849 53359
rect 60895 53313 60973 53359
rect 61019 53313 61097 53359
rect 61143 53313 61221 53359
rect 61267 53313 61345 53359
rect 61391 53313 61469 53359
rect 61515 53313 61593 53359
rect 61639 53313 61717 53359
rect 61763 53313 61841 53359
rect 61887 53313 61965 53359
rect 62011 53313 62089 53359
rect 62135 53313 62213 53359
rect 62259 53313 62337 53359
rect 62383 53313 62461 53359
rect 62507 53313 62585 53359
rect 62631 53313 62709 53359
rect 62755 53313 62833 53359
rect 62879 53313 62957 53359
rect 63003 53313 63081 53359
rect 63127 53313 63205 53359
rect 63251 53313 63329 53359
rect 63375 53313 63453 53359
rect 63499 53313 63577 53359
rect 63623 53313 63701 53359
rect 63747 53313 63825 53359
rect 63871 53313 63949 53359
rect 63995 53313 64073 53359
rect 64119 53313 64197 53359
rect 64243 53313 64321 53359
rect 64367 53313 64445 53359
rect 64491 53313 64569 53359
rect 64615 53313 64693 53359
rect 64739 53313 64817 53359
rect 64863 53313 64941 53359
rect 64987 53313 65065 53359
rect 65111 53313 65189 53359
rect 65235 53313 65313 53359
rect 65359 53313 65437 53359
rect 65483 53313 65561 53359
rect 65607 53313 65685 53359
rect 65731 53313 65809 53359
rect 65855 53313 65933 53359
rect 65979 53313 66057 53359
rect 66103 53313 66181 53359
rect 66227 53313 66305 53359
rect 66351 53313 66429 53359
rect 66475 53313 66553 53359
rect 66599 53313 66677 53359
rect 66723 53313 66801 53359
rect 66847 53313 66925 53359
rect 66971 53313 67049 53359
rect 67095 53313 67173 53359
rect 67219 53313 67297 53359
rect 67343 53313 67421 53359
rect 67467 53313 67545 53359
rect 67591 53313 67669 53359
rect 67715 53313 67793 53359
rect 67839 53313 67917 53359
rect 67963 53313 68041 53359
rect 68087 53313 68165 53359
rect 68211 53313 68289 53359
rect 68335 53313 68413 53359
rect 68459 53313 68537 53359
rect 68583 53313 68661 53359
rect 68707 53313 68785 53359
rect 68831 53313 68909 53359
rect 68955 53313 69033 53359
rect 69079 53313 69157 53359
rect 69203 53313 69281 53359
rect 69327 53313 69405 53359
rect 69451 53313 69529 53359
rect 69575 53313 69653 53359
rect 69699 53313 69777 53359
rect 69823 53313 69901 53359
rect 69947 53313 70025 53359
rect 70071 53313 70149 53359
rect 70195 53313 70273 53359
rect 70319 53313 70397 53359
rect 70443 53313 70521 53359
rect 70567 53313 70645 53359
rect 70691 53313 70769 53359
rect 70815 53313 70893 53359
rect 70939 53313 71017 53359
rect 71063 53313 71141 53359
rect 71187 53313 71265 53359
rect 71311 53313 71389 53359
rect 71435 53313 71513 53359
rect 71559 53313 71637 53359
rect 71683 53313 71761 53359
rect 71807 53313 71885 53359
rect 71931 53313 72009 53359
rect 72055 53313 72133 53359
rect 72179 53313 72257 53359
rect 72303 53313 72381 53359
rect 72427 53313 72505 53359
rect 72551 53313 72629 53359
rect 72675 53313 72753 53359
rect 72799 53313 72877 53359
rect 72923 53313 73001 53359
rect 73047 53313 73125 53359
rect 73171 53313 73249 53359
rect 73295 53313 73373 53359
rect 73419 53313 73497 53359
rect 73543 53313 73621 53359
rect 73667 53313 73745 53359
rect 73791 53313 73869 53359
rect 73915 53313 73993 53359
rect 74039 53313 74117 53359
rect 74163 53313 74241 53359
rect 74287 53313 74365 53359
rect 74411 53313 74489 53359
rect 74535 53313 74613 53359
rect 74659 53313 74737 53359
rect 74783 53313 74861 53359
rect 74907 53313 74985 53359
rect 75031 53313 75109 53359
rect 75155 53313 75233 53359
rect 75279 53313 75357 53359
rect 75403 53313 75481 53359
rect 75527 53313 75605 53359
rect 75651 53313 75729 53359
rect 75775 53313 75853 53359
rect 75899 53313 75977 53359
rect 76023 53313 76101 53359
rect 76147 53313 76225 53359
rect 76271 53313 76349 53359
rect 76395 53313 76473 53359
rect 76519 53313 76597 53359
rect 76643 53313 76721 53359
rect 76767 53313 76845 53359
rect 76891 53313 76969 53359
rect 77015 53313 77093 53359
rect 77139 53313 77217 53359
rect 77263 53313 77341 53359
rect 77387 53313 77465 53359
rect 77511 53313 77589 53359
rect 77635 53313 77713 53359
rect 77759 53313 77837 53359
rect 77883 53313 77961 53359
rect 78007 53313 78085 53359
rect 78131 53313 78209 53359
rect 78255 53313 78333 53359
rect 78379 53313 78457 53359
rect 78503 53313 78581 53359
rect 78627 53313 78705 53359
rect 78751 53313 78829 53359
rect 78875 53313 78953 53359
rect 78999 53313 79077 53359
rect 79123 53313 79201 53359
rect 79247 53313 79325 53359
rect 79371 53313 79449 53359
rect 79495 53313 79573 53359
rect 79619 53313 79697 53359
rect 79743 53313 79821 53359
rect 79867 53313 79945 53359
rect 79991 53313 80069 53359
rect 80115 53313 80193 53359
rect 80239 53313 80317 53359
rect 80363 53313 80441 53359
rect 80487 53313 80565 53359
rect 80611 53313 80689 53359
rect 80735 53313 80813 53359
rect 80859 53313 80937 53359
rect 80983 53313 81061 53359
rect 81107 53313 81185 53359
rect 81231 53313 81309 53359
rect 81355 53313 81433 53359
rect 81479 53313 81557 53359
rect 81603 53313 81681 53359
rect 81727 53313 81805 53359
rect 81851 53313 81929 53359
rect 81975 53313 82053 53359
rect 82099 53313 82177 53359
rect 82223 53313 82301 53359
rect 82347 53313 82425 53359
rect 82471 53313 82549 53359
rect 82595 53313 82673 53359
rect 82719 53313 82797 53359
rect 82843 53313 82921 53359
rect 82967 53313 83045 53359
rect 83091 53313 83169 53359
rect 83215 53313 83293 53359
rect 83339 53313 83417 53359
rect 83463 53313 83541 53359
rect 83587 53313 83665 53359
rect 83711 53313 83789 53359
rect 83835 53313 83913 53359
rect 83959 53313 84037 53359
rect 84083 53313 84161 53359
rect 84207 53313 84285 53359
rect 84331 53313 84409 53359
rect 84455 53313 84533 53359
rect 84579 53313 84657 53359
rect 84703 53313 84781 53359
rect 84827 53313 84905 53359
rect 84951 53313 85029 53359
rect 85075 53313 85153 53359
rect 85199 53313 85277 53359
rect 85323 53313 85401 53359
rect 85447 53313 85525 53359
rect 85571 53313 85649 53359
rect 85695 53313 85816 53359
rect 70 53235 85816 53313
rect 70 53189 89 53235
rect 135 53189 213 53235
rect 259 53189 337 53235
rect 383 53189 461 53235
rect 507 53189 585 53235
rect 631 53189 709 53235
rect 755 53189 833 53235
rect 879 53189 957 53235
rect 1003 53189 1081 53235
rect 1127 53189 1205 53235
rect 1251 53189 1329 53235
rect 1375 53189 1453 53235
rect 1499 53189 1577 53235
rect 1623 53189 1701 53235
rect 1747 53189 1825 53235
rect 1871 53189 1949 53235
rect 1995 53189 2073 53235
rect 2119 53189 2197 53235
rect 2243 53189 2321 53235
rect 2367 53189 2445 53235
rect 2491 53189 2569 53235
rect 2615 53189 2693 53235
rect 2739 53189 2817 53235
rect 2863 53189 2941 53235
rect 2987 53189 3065 53235
rect 3111 53189 3189 53235
rect 3235 53189 3313 53235
rect 3359 53189 3437 53235
rect 3483 53189 3561 53235
rect 3607 53189 3685 53235
rect 3731 53189 3809 53235
rect 3855 53189 3933 53235
rect 3979 53189 4057 53235
rect 4103 53189 4181 53235
rect 4227 53189 4305 53235
rect 4351 53189 4429 53235
rect 4475 53189 4553 53235
rect 4599 53189 4677 53235
rect 4723 53189 4801 53235
rect 4847 53189 4925 53235
rect 4971 53189 5049 53235
rect 5095 53189 5173 53235
rect 5219 53189 5297 53235
rect 5343 53189 5421 53235
rect 5467 53189 5545 53235
rect 5591 53189 5669 53235
rect 5715 53189 5793 53235
rect 5839 53189 5917 53235
rect 5963 53189 6041 53235
rect 6087 53189 6165 53235
rect 6211 53189 6289 53235
rect 6335 53189 6413 53235
rect 6459 53189 6537 53235
rect 6583 53189 6661 53235
rect 6707 53189 6785 53235
rect 6831 53189 6909 53235
rect 6955 53189 7033 53235
rect 7079 53189 7157 53235
rect 7203 53189 7281 53235
rect 7327 53189 7405 53235
rect 7451 53189 7529 53235
rect 7575 53189 7653 53235
rect 7699 53189 7777 53235
rect 7823 53189 7901 53235
rect 7947 53189 8025 53235
rect 8071 53189 8149 53235
rect 8195 53189 8273 53235
rect 8319 53189 8397 53235
rect 8443 53189 8521 53235
rect 8567 53189 8645 53235
rect 8691 53189 8769 53235
rect 8815 53189 8893 53235
rect 8939 53189 9017 53235
rect 9063 53189 9141 53235
rect 9187 53189 9265 53235
rect 9311 53189 9389 53235
rect 9435 53189 9513 53235
rect 9559 53189 9637 53235
rect 9683 53189 9761 53235
rect 9807 53189 9885 53235
rect 9931 53189 10009 53235
rect 10055 53189 10133 53235
rect 10179 53189 10257 53235
rect 10303 53189 10381 53235
rect 10427 53189 10505 53235
rect 10551 53189 10629 53235
rect 10675 53189 10753 53235
rect 10799 53189 10877 53235
rect 10923 53189 11001 53235
rect 11047 53189 11125 53235
rect 11171 53189 11249 53235
rect 11295 53189 11373 53235
rect 11419 53189 11497 53235
rect 11543 53189 11621 53235
rect 11667 53189 11745 53235
rect 11791 53189 11869 53235
rect 11915 53189 11993 53235
rect 12039 53189 12117 53235
rect 12163 53189 12241 53235
rect 12287 53189 12365 53235
rect 12411 53189 12489 53235
rect 12535 53189 12613 53235
rect 12659 53189 12737 53235
rect 12783 53189 12861 53235
rect 12907 53189 12985 53235
rect 13031 53189 13109 53235
rect 13155 53189 13233 53235
rect 13279 53189 13357 53235
rect 13403 53189 13481 53235
rect 13527 53189 13605 53235
rect 13651 53189 13729 53235
rect 13775 53189 13853 53235
rect 13899 53189 13977 53235
rect 14023 53189 14101 53235
rect 14147 53189 14225 53235
rect 14271 53189 14349 53235
rect 14395 53189 14473 53235
rect 14519 53189 14597 53235
rect 14643 53189 14721 53235
rect 14767 53189 14845 53235
rect 14891 53189 14969 53235
rect 15015 53189 15093 53235
rect 15139 53189 15217 53235
rect 15263 53189 15341 53235
rect 15387 53189 15465 53235
rect 15511 53189 15589 53235
rect 15635 53189 15713 53235
rect 15759 53189 15837 53235
rect 15883 53189 15961 53235
rect 16007 53189 16085 53235
rect 16131 53189 16209 53235
rect 16255 53189 16333 53235
rect 16379 53189 16457 53235
rect 16503 53189 16581 53235
rect 16627 53189 16705 53235
rect 16751 53189 16829 53235
rect 16875 53189 16953 53235
rect 16999 53189 17077 53235
rect 17123 53189 17201 53235
rect 17247 53189 17325 53235
rect 17371 53189 17449 53235
rect 17495 53189 17573 53235
rect 17619 53189 17697 53235
rect 17743 53189 17821 53235
rect 17867 53189 17945 53235
rect 17991 53189 18069 53235
rect 18115 53189 18193 53235
rect 18239 53189 18317 53235
rect 18363 53189 18441 53235
rect 18487 53189 18565 53235
rect 18611 53189 18689 53235
rect 18735 53189 18813 53235
rect 18859 53189 18937 53235
rect 18983 53189 19061 53235
rect 19107 53189 19185 53235
rect 19231 53189 19309 53235
rect 19355 53189 19433 53235
rect 19479 53189 19557 53235
rect 19603 53189 19681 53235
rect 19727 53189 19805 53235
rect 19851 53189 19929 53235
rect 19975 53189 20053 53235
rect 20099 53189 20177 53235
rect 20223 53189 20301 53235
rect 20347 53189 20425 53235
rect 20471 53189 20549 53235
rect 20595 53189 20673 53235
rect 20719 53189 20797 53235
rect 20843 53189 20921 53235
rect 20967 53189 21045 53235
rect 21091 53189 21169 53235
rect 21215 53189 21293 53235
rect 21339 53189 21417 53235
rect 21463 53189 21541 53235
rect 21587 53189 21665 53235
rect 21711 53189 21789 53235
rect 21835 53189 21913 53235
rect 21959 53189 22037 53235
rect 22083 53189 22161 53235
rect 22207 53189 22285 53235
rect 22331 53189 22409 53235
rect 22455 53189 22533 53235
rect 22579 53189 22657 53235
rect 22703 53189 22781 53235
rect 22827 53189 22905 53235
rect 22951 53189 23029 53235
rect 23075 53189 23153 53235
rect 23199 53189 23277 53235
rect 23323 53189 23401 53235
rect 23447 53189 23525 53235
rect 23571 53189 23649 53235
rect 23695 53189 23773 53235
rect 23819 53189 23897 53235
rect 23943 53189 24021 53235
rect 24067 53189 24145 53235
rect 24191 53189 24269 53235
rect 24315 53189 24393 53235
rect 24439 53189 24517 53235
rect 24563 53189 24641 53235
rect 24687 53189 24765 53235
rect 24811 53189 24889 53235
rect 24935 53189 25013 53235
rect 25059 53189 25137 53235
rect 25183 53189 25261 53235
rect 25307 53189 25385 53235
rect 25431 53189 25509 53235
rect 25555 53189 25633 53235
rect 25679 53189 25757 53235
rect 25803 53189 25881 53235
rect 25927 53189 26005 53235
rect 26051 53189 26129 53235
rect 26175 53189 26253 53235
rect 26299 53189 26377 53235
rect 26423 53189 26501 53235
rect 26547 53189 26625 53235
rect 26671 53189 26749 53235
rect 26795 53189 26873 53235
rect 26919 53189 26997 53235
rect 27043 53189 27121 53235
rect 27167 53189 27245 53235
rect 27291 53189 27369 53235
rect 27415 53189 27493 53235
rect 27539 53189 27617 53235
rect 27663 53189 27741 53235
rect 27787 53189 27865 53235
rect 27911 53189 27989 53235
rect 28035 53189 28113 53235
rect 28159 53189 28237 53235
rect 28283 53189 28361 53235
rect 28407 53189 28485 53235
rect 28531 53189 28609 53235
rect 28655 53189 28733 53235
rect 28779 53189 28857 53235
rect 28903 53189 28981 53235
rect 29027 53189 29105 53235
rect 29151 53189 29229 53235
rect 29275 53189 29353 53235
rect 29399 53189 29477 53235
rect 29523 53189 29601 53235
rect 29647 53189 29725 53235
rect 29771 53189 29849 53235
rect 29895 53189 29973 53235
rect 30019 53189 30097 53235
rect 30143 53189 30221 53235
rect 30267 53189 30345 53235
rect 30391 53189 30469 53235
rect 30515 53189 30593 53235
rect 30639 53189 30717 53235
rect 30763 53189 30841 53235
rect 30887 53189 30965 53235
rect 31011 53189 31089 53235
rect 31135 53189 31213 53235
rect 31259 53189 31337 53235
rect 31383 53189 31461 53235
rect 31507 53189 31585 53235
rect 31631 53189 31709 53235
rect 31755 53189 31833 53235
rect 31879 53189 31957 53235
rect 32003 53189 32081 53235
rect 32127 53189 32205 53235
rect 32251 53189 32329 53235
rect 32375 53189 32453 53235
rect 32499 53189 32577 53235
rect 32623 53189 32701 53235
rect 32747 53189 32825 53235
rect 32871 53189 32949 53235
rect 32995 53189 33073 53235
rect 33119 53189 33197 53235
rect 33243 53189 33321 53235
rect 33367 53189 33445 53235
rect 33491 53189 33569 53235
rect 33615 53189 33693 53235
rect 33739 53189 33817 53235
rect 33863 53189 33941 53235
rect 33987 53189 34065 53235
rect 34111 53189 34189 53235
rect 34235 53189 34313 53235
rect 34359 53189 34437 53235
rect 34483 53189 34561 53235
rect 34607 53189 34685 53235
rect 34731 53189 34809 53235
rect 34855 53189 34933 53235
rect 34979 53189 35057 53235
rect 35103 53189 35181 53235
rect 35227 53189 35305 53235
rect 35351 53189 35429 53235
rect 35475 53189 35553 53235
rect 35599 53189 35677 53235
rect 35723 53189 35801 53235
rect 35847 53189 35925 53235
rect 35971 53189 36049 53235
rect 36095 53189 36173 53235
rect 36219 53189 36297 53235
rect 36343 53189 36421 53235
rect 36467 53189 36545 53235
rect 36591 53189 36669 53235
rect 36715 53189 36793 53235
rect 36839 53189 36917 53235
rect 36963 53189 37041 53235
rect 37087 53189 37165 53235
rect 37211 53189 37289 53235
rect 37335 53189 37413 53235
rect 37459 53189 37537 53235
rect 37583 53189 37661 53235
rect 37707 53189 37785 53235
rect 37831 53189 37909 53235
rect 37955 53189 38033 53235
rect 38079 53189 38157 53235
rect 38203 53189 38281 53235
rect 38327 53189 38405 53235
rect 38451 53189 38529 53235
rect 38575 53189 38653 53235
rect 38699 53189 38777 53235
rect 38823 53189 38901 53235
rect 38947 53189 39025 53235
rect 39071 53189 39149 53235
rect 39195 53189 39273 53235
rect 39319 53189 39397 53235
rect 39443 53189 39521 53235
rect 39567 53189 39645 53235
rect 39691 53189 39769 53235
rect 39815 53189 39893 53235
rect 39939 53189 40017 53235
rect 40063 53189 40141 53235
rect 40187 53189 40265 53235
rect 40311 53189 40389 53235
rect 40435 53189 40513 53235
rect 40559 53189 40637 53235
rect 40683 53189 40761 53235
rect 40807 53189 40885 53235
rect 40931 53189 41009 53235
rect 41055 53189 41133 53235
rect 41179 53189 41257 53235
rect 41303 53189 41381 53235
rect 41427 53189 41505 53235
rect 41551 53189 41629 53235
rect 41675 53189 41753 53235
rect 41799 53189 41877 53235
rect 41923 53189 42001 53235
rect 42047 53189 42125 53235
rect 42171 53189 42249 53235
rect 42295 53189 42373 53235
rect 42419 53189 42497 53235
rect 42543 53189 42621 53235
rect 42667 53189 42745 53235
rect 42791 53189 42869 53235
rect 42915 53189 42993 53235
rect 43039 53189 43117 53235
rect 43163 53189 43241 53235
rect 43287 53189 43365 53235
rect 43411 53189 43489 53235
rect 43535 53189 43613 53235
rect 43659 53189 43737 53235
rect 43783 53189 43861 53235
rect 43907 53189 43985 53235
rect 44031 53189 44109 53235
rect 44155 53189 44233 53235
rect 44279 53189 44357 53235
rect 44403 53189 44481 53235
rect 44527 53189 44605 53235
rect 44651 53189 44729 53235
rect 44775 53189 44853 53235
rect 44899 53189 44977 53235
rect 45023 53189 45101 53235
rect 45147 53189 45225 53235
rect 45271 53189 45349 53235
rect 45395 53189 45473 53235
rect 45519 53189 45597 53235
rect 45643 53189 45721 53235
rect 45767 53189 45845 53235
rect 45891 53189 45969 53235
rect 46015 53189 46093 53235
rect 46139 53189 46217 53235
rect 46263 53189 46341 53235
rect 46387 53189 46465 53235
rect 46511 53189 46589 53235
rect 46635 53189 46713 53235
rect 46759 53189 46837 53235
rect 46883 53189 46961 53235
rect 47007 53189 47085 53235
rect 47131 53189 47209 53235
rect 47255 53189 47333 53235
rect 47379 53189 47457 53235
rect 47503 53189 47581 53235
rect 47627 53189 47705 53235
rect 47751 53189 47829 53235
rect 47875 53189 47953 53235
rect 47999 53189 48077 53235
rect 48123 53189 48201 53235
rect 48247 53189 48325 53235
rect 48371 53189 48449 53235
rect 48495 53189 48573 53235
rect 48619 53189 48697 53235
rect 48743 53189 48821 53235
rect 48867 53189 48945 53235
rect 48991 53189 49069 53235
rect 49115 53189 49193 53235
rect 49239 53189 49317 53235
rect 49363 53189 49441 53235
rect 49487 53189 49565 53235
rect 49611 53189 49689 53235
rect 49735 53189 49813 53235
rect 49859 53189 49937 53235
rect 49983 53189 50061 53235
rect 50107 53189 50185 53235
rect 50231 53189 50309 53235
rect 50355 53189 50433 53235
rect 50479 53189 50557 53235
rect 50603 53189 50681 53235
rect 50727 53189 50805 53235
rect 50851 53189 50929 53235
rect 50975 53189 51053 53235
rect 51099 53189 51177 53235
rect 51223 53189 51301 53235
rect 51347 53189 51425 53235
rect 51471 53189 51549 53235
rect 51595 53189 51673 53235
rect 51719 53189 51797 53235
rect 51843 53189 51921 53235
rect 51967 53189 52045 53235
rect 52091 53189 52169 53235
rect 52215 53189 52293 53235
rect 52339 53189 52417 53235
rect 52463 53189 52541 53235
rect 52587 53189 52665 53235
rect 52711 53189 52789 53235
rect 52835 53189 52913 53235
rect 52959 53189 53037 53235
rect 53083 53189 53161 53235
rect 53207 53189 53285 53235
rect 53331 53189 53409 53235
rect 53455 53189 53533 53235
rect 53579 53189 53657 53235
rect 53703 53189 53781 53235
rect 53827 53189 53905 53235
rect 53951 53189 54029 53235
rect 54075 53189 54153 53235
rect 54199 53189 54277 53235
rect 54323 53189 54401 53235
rect 54447 53189 54525 53235
rect 54571 53189 54649 53235
rect 54695 53189 54773 53235
rect 54819 53189 54897 53235
rect 54943 53189 55021 53235
rect 55067 53189 55145 53235
rect 55191 53189 55269 53235
rect 55315 53189 55393 53235
rect 55439 53189 55517 53235
rect 55563 53189 55641 53235
rect 55687 53189 55765 53235
rect 55811 53189 55889 53235
rect 55935 53189 56013 53235
rect 56059 53189 56137 53235
rect 56183 53189 56261 53235
rect 56307 53189 56385 53235
rect 56431 53189 56509 53235
rect 56555 53189 56633 53235
rect 56679 53189 56757 53235
rect 56803 53189 56881 53235
rect 56927 53189 57005 53235
rect 57051 53189 57129 53235
rect 57175 53189 57253 53235
rect 57299 53189 57377 53235
rect 57423 53189 57501 53235
rect 57547 53189 57625 53235
rect 57671 53189 57749 53235
rect 57795 53189 57873 53235
rect 57919 53189 57997 53235
rect 58043 53189 58121 53235
rect 58167 53189 58245 53235
rect 58291 53189 58369 53235
rect 58415 53189 58493 53235
rect 58539 53189 58617 53235
rect 58663 53189 58741 53235
rect 58787 53189 58865 53235
rect 58911 53189 58989 53235
rect 59035 53189 59113 53235
rect 59159 53189 59237 53235
rect 59283 53189 59361 53235
rect 59407 53189 59485 53235
rect 59531 53189 59609 53235
rect 59655 53189 59733 53235
rect 59779 53189 59857 53235
rect 59903 53189 59981 53235
rect 60027 53189 60105 53235
rect 60151 53189 60229 53235
rect 60275 53189 60353 53235
rect 60399 53189 60477 53235
rect 60523 53189 60601 53235
rect 60647 53189 60725 53235
rect 60771 53189 60849 53235
rect 60895 53189 60973 53235
rect 61019 53189 61097 53235
rect 61143 53189 61221 53235
rect 61267 53189 61345 53235
rect 61391 53189 61469 53235
rect 61515 53189 61593 53235
rect 61639 53189 61717 53235
rect 61763 53189 61841 53235
rect 61887 53189 61965 53235
rect 62011 53189 62089 53235
rect 62135 53189 62213 53235
rect 62259 53189 62337 53235
rect 62383 53189 62461 53235
rect 62507 53189 62585 53235
rect 62631 53189 62709 53235
rect 62755 53189 62833 53235
rect 62879 53189 62957 53235
rect 63003 53189 63081 53235
rect 63127 53189 63205 53235
rect 63251 53189 63329 53235
rect 63375 53189 63453 53235
rect 63499 53189 63577 53235
rect 63623 53189 63701 53235
rect 63747 53189 63825 53235
rect 63871 53189 63949 53235
rect 63995 53189 64073 53235
rect 64119 53189 64197 53235
rect 64243 53189 64321 53235
rect 64367 53189 64445 53235
rect 64491 53189 64569 53235
rect 64615 53189 64693 53235
rect 64739 53189 64817 53235
rect 64863 53189 64941 53235
rect 64987 53189 65065 53235
rect 65111 53189 65189 53235
rect 65235 53189 65313 53235
rect 65359 53189 65437 53235
rect 65483 53189 65561 53235
rect 65607 53189 65685 53235
rect 65731 53189 65809 53235
rect 65855 53189 65933 53235
rect 65979 53189 66057 53235
rect 66103 53189 66181 53235
rect 66227 53189 66305 53235
rect 66351 53189 66429 53235
rect 66475 53189 66553 53235
rect 66599 53189 66677 53235
rect 66723 53189 66801 53235
rect 66847 53189 66925 53235
rect 66971 53189 67049 53235
rect 67095 53189 67173 53235
rect 67219 53189 67297 53235
rect 67343 53189 67421 53235
rect 67467 53189 67545 53235
rect 67591 53189 67669 53235
rect 67715 53189 67793 53235
rect 67839 53189 67917 53235
rect 67963 53189 68041 53235
rect 68087 53189 68165 53235
rect 68211 53189 68289 53235
rect 68335 53189 68413 53235
rect 68459 53189 68537 53235
rect 68583 53189 68661 53235
rect 68707 53189 68785 53235
rect 68831 53189 68909 53235
rect 68955 53189 69033 53235
rect 69079 53189 69157 53235
rect 69203 53189 69281 53235
rect 69327 53189 69405 53235
rect 69451 53189 69529 53235
rect 69575 53189 69653 53235
rect 69699 53189 69777 53235
rect 69823 53189 69901 53235
rect 69947 53189 70025 53235
rect 70071 53189 70149 53235
rect 70195 53189 70273 53235
rect 70319 53189 70397 53235
rect 70443 53189 70521 53235
rect 70567 53189 70645 53235
rect 70691 53189 70769 53235
rect 70815 53189 70893 53235
rect 70939 53189 71017 53235
rect 71063 53189 71141 53235
rect 71187 53189 71265 53235
rect 71311 53189 71389 53235
rect 71435 53189 71513 53235
rect 71559 53189 71637 53235
rect 71683 53189 71761 53235
rect 71807 53189 71885 53235
rect 71931 53189 72009 53235
rect 72055 53189 72133 53235
rect 72179 53189 72257 53235
rect 72303 53189 72381 53235
rect 72427 53189 72505 53235
rect 72551 53189 72629 53235
rect 72675 53189 72753 53235
rect 72799 53189 72877 53235
rect 72923 53189 73001 53235
rect 73047 53189 73125 53235
rect 73171 53189 73249 53235
rect 73295 53189 73373 53235
rect 73419 53189 73497 53235
rect 73543 53189 73621 53235
rect 73667 53189 73745 53235
rect 73791 53189 73869 53235
rect 73915 53189 73993 53235
rect 74039 53189 74117 53235
rect 74163 53189 74241 53235
rect 74287 53189 74365 53235
rect 74411 53189 74489 53235
rect 74535 53189 74613 53235
rect 74659 53189 74737 53235
rect 74783 53189 74861 53235
rect 74907 53189 74985 53235
rect 75031 53189 75109 53235
rect 75155 53189 75233 53235
rect 75279 53189 75357 53235
rect 75403 53189 75481 53235
rect 75527 53189 75605 53235
rect 75651 53189 75729 53235
rect 75775 53189 75853 53235
rect 75899 53189 75977 53235
rect 76023 53189 76101 53235
rect 76147 53189 76225 53235
rect 76271 53189 76349 53235
rect 76395 53189 76473 53235
rect 76519 53189 76597 53235
rect 76643 53189 76721 53235
rect 76767 53189 76845 53235
rect 76891 53189 76969 53235
rect 77015 53189 77093 53235
rect 77139 53189 77217 53235
rect 77263 53189 77341 53235
rect 77387 53189 77465 53235
rect 77511 53189 77589 53235
rect 77635 53189 77713 53235
rect 77759 53189 77837 53235
rect 77883 53189 77961 53235
rect 78007 53189 78085 53235
rect 78131 53189 78209 53235
rect 78255 53189 78333 53235
rect 78379 53189 78457 53235
rect 78503 53189 78581 53235
rect 78627 53189 78705 53235
rect 78751 53189 78829 53235
rect 78875 53189 78953 53235
rect 78999 53189 79077 53235
rect 79123 53189 79201 53235
rect 79247 53189 79325 53235
rect 79371 53189 79449 53235
rect 79495 53189 79573 53235
rect 79619 53189 79697 53235
rect 79743 53189 79821 53235
rect 79867 53189 79945 53235
rect 79991 53189 80069 53235
rect 80115 53189 80193 53235
rect 80239 53189 80317 53235
rect 80363 53189 80441 53235
rect 80487 53189 80565 53235
rect 80611 53189 80689 53235
rect 80735 53189 80813 53235
rect 80859 53189 80937 53235
rect 80983 53189 81061 53235
rect 81107 53189 81185 53235
rect 81231 53189 81309 53235
rect 81355 53189 81433 53235
rect 81479 53189 81557 53235
rect 81603 53189 81681 53235
rect 81727 53189 81805 53235
rect 81851 53189 81929 53235
rect 81975 53189 82053 53235
rect 82099 53189 82177 53235
rect 82223 53189 82301 53235
rect 82347 53189 82425 53235
rect 82471 53189 82549 53235
rect 82595 53189 82673 53235
rect 82719 53189 82797 53235
rect 82843 53189 82921 53235
rect 82967 53189 83045 53235
rect 83091 53189 83169 53235
rect 83215 53189 83293 53235
rect 83339 53189 83417 53235
rect 83463 53189 83541 53235
rect 83587 53189 83665 53235
rect 83711 53189 83789 53235
rect 83835 53189 83913 53235
rect 83959 53189 84037 53235
rect 84083 53189 84161 53235
rect 84207 53189 84285 53235
rect 84331 53189 84409 53235
rect 84455 53189 84533 53235
rect 84579 53189 84657 53235
rect 84703 53189 84781 53235
rect 84827 53189 84905 53235
rect 84951 53189 85029 53235
rect 85075 53189 85153 53235
rect 85199 53189 85277 53235
rect 85323 53189 85401 53235
rect 85447 53189 85525 53235
rect 85571 53189 85649 53235
rect 85695 53189 85816 53235
rect 70 53111 85816 53189
rect 70 53065 89 53111
rect 135 53065 213 53111
rect 259 53065 337 53111
rect 383 53065 461 53111
rect 507 53065 585 53111
rect 631 53065 709 53111
rect 755 53065 833 53111
rect 879 53065 957 53111
rect 1003 53065 1081 53111
rect 1127 53065 1205 53111
rect 1251 53065 1329 53111
rect 1375 53065 1453 53111
rect 1499 53065 1577 53111
rect 1623 53065 1701 53111
rect 1747 53065 1825 53111
rect 1871 53065 1949 53111
rect 1995 53065 2073 53111
rect 2119 53065 2197 53111
rect 2243 53065 2321 53111
rect 2367 53065 2445 53111
rect 2491 53065 2569 53111
rect 2615 53065 2693 53111
rect 2739 53065 2817 53111
rect 2863 53065 2941 53111
rect 2987 53065 3065 53111
rect 3111 53065 3189 53111
rect 3235 53065 3313 53111
rect 3359 53065 3437 53111
rect 3483 53065 3561 53111
rect 3607 53065 3685 53111
rect 3731 53065 3809 53111
rect 3855 53065 3933 53111
rect 3979 53065 4057 53111
rect 4103 53065 4181 53111
rect 4227 53065 4305 53111
rect 4351 53065 4429 53111
rect 4475 53065 4553 53111
rect 4599 53065 4677 53111
rect 4723 53065 4801 53111
rect 4847 53065 4925 53111
rect 4971 53065 5049 53111
rect 5095 53065 5173 53111
rect 5219 53065 5297 53111
rect 5343 53065 5421 53111
rect 5467 53065 5545 53111
rect 5591 53065 5669 53111
rect 5715 53065 5793 53111
rect 5839 53065 5917 53111
rect 5963 53065 6041 53111
rect 6087 53065 6165 53111
rect 6211 53065 6289 53111
rect 6335 53065 6413 53111
rect 6459 53065 6537 53111
rect 6583 53065 6661 53111
rect 6707 53065 6785 53111
rect 6831 53065 6909 53111
rect 6955 53065 7033 53111
rect 7079 53065 7157 53111
rect 7203 53065 7281 53111
rect 7327 53065 7405 53111
rect 7451 53065 7529 53111
rect 7575 53065 7653 53111
rect 7699 53065 7777 53111
rect 7823 53065 7901 53111
rect 7947 53065 8025 53111
rect 8071 53065 8149 53111
rect 8195 53065 8273 53111
rect 8319 53065 8397 53111
rect 8443 53065 8521 53111
rect 8567 53065 8645 53111
rect 8691 53065 8769 53111
rect 8815 53065 8893 53111
rect 8939 53065 9017 53111
rect 9063 53065 9141 53111
rect 9187 53065 9265 53111
rect 9311 53065 9389 53111
rect 9435 53065 9513 53111
rect 9559 53065 9637 53111
rect 9683 53065 9761 53111
rect 9807 53065 9885 53111
rect 9931 53065 10009 53111
rect 10055 53065 10133 53111
rect 10179 53065 10257 53111
rect 10303 53065 10381 53111
rect 10427 53065 10505 53111
rect 10551 53065 10629 53111
rect 10675 53065 10753 53111
rect 10799 53065 10877 53111
rect 10923 53065 11001 53111
rect 11047 53065 11125 53111
rect 11171 53065 11249 53111
rect 11295 53065 11373 53111
rect 11419 53065 11497 53111
rect 11543 53065 11621 53111
rect 11667 53065 11745 53111
rect 11791 53065 11869 53111
rect 11915 53065 11993 53111
rect 12039 53065 12117 53111
rect 12163 53065 12241 53111
rect 12287 53065 12365 53111
rect 12411 53065 12489 53111
rect 12535 53065 12613 53111
rect 12659 53065 12737 53111
rect 12783 53065 12861 53111
rect 12907 53065 12985 53111
rect 13031 53065 13109 53111
rect 13155 53065 13233 53111
rect 13279 53065 13357 53111
rect 13403 53065 13481 53111
rect 13527 53065 13605 53111
rect 13651 53065 13729 53111
rect 13775 53065 13853 53111
rect 13899 53065 13977 53111
rect 14023 53065 14101 53111
rect 14147 53065 14225 53111
rect 14271 53065 14349 53111
rect 14395 53065 14473 53111
rect 14519 53065 14597 53111
rect 14643 53065 14721 53111
rect 14767 53065 14845 53111
rect 14891 53065 14969 53111
rect 15015 53065 15093 53111
rect 15139 53065 15217 53111
rect 15263 53065 15341 53111
rect 15387 53065 15465 53111
rect 15511 53065 15589 53111
rect 15635 53065 15713 53111
rect 15759 53065 15837 53111
rect 15883 53065 15961 53111
rect 16007 53065 16085 53111
rect 16131 53065 16209 53111
rect 16255 53065 16333 53111
rect 16379 53065 16457 53111
rect 16503 53065 16581 53111
rect 16627 53065 16705 53111
rect 16751 53065 16829 53111
rect 16875 53065 16953 53111
rect 16999 53065 17077 53111
rect 17123 53065 17201 53111
rect 17247 53065 17325 53111
rect 17371 53065 17449 53111
rect 17495 53065 17573 53111
rect 17619 53065 17697 53111
rect 17743 53065 17821 53111
rect 17867 53065 17945 53111
rect 17991 53065 18069 53111
rect 18115 53065 18193 53111
rect 18239 53065 18317 53111
rect 18363 53065 18441 53111
rect 18487 53065 18565 53111
rect 18611 53065 18689 53111
rect 18735 53065 18813 53111
rect 18859 53065 18937 53111
rect 18983 53065 19061 53111
rect 19107 53065 19185 53111
rect 19231 53065 19309 53111
rect 19355 53065 19433 53111
rect 19479 53065 19557 53111
rect 19603 53065 19681 53111
rect 19727 53065 19805 53111
rect 19851 53065 19929 53111
rect 19975 53065 20053 53111
rect 20099 53065 20177 53111
rect 20223 53065 20301 53111
rect 20347 53065 20425 53111
rect 20471 53065 20549 53111
rect 20595 53065 20673 53111
rect 20719 53065 20797 53111
rect 20843 53065 20921 53111
rect 20967 53065 21045 53111
rect 21091 53065 21169 53111
rect 21215 53065 21293 53111
rect 21339 53065 21417 53111
rect 21463 53065 21541 53111
rect 21587 53065 21665 53111
rect 21711 53065 21789 53111
rect 21835 53065 21913 53111
rect 21959 53065 22037 53111
rect 22083 53065 22161 53111
rect 22207 53065 22285 53111
rect 22331 53065 22409 53111
rect 22455 53065 22533 53111
rect 22579 53065 22657 53111
rect 22703 53065 22781 53111
rect 22827 53065 22905 53111
rect 22951 53065 23029 53111
rect 23075 53065 23153 53111
rect 23199 53065 23277 53111
rect 23323 53065 23401 53111
rect 23447 53065 23525 53111
rect 23571 53065 23649 53111
rect 23695 53065 23773 53111
rect 23819 53065 23897 53111
rect 23943 53065 24021 53111
rect 24067 53065 24145 53111
rect 24191 53065 24269 53111
rect 24315 53065 24393 53111
rect 24439 53065 24517 53111
rect 24563 53065 24641 53111
rect 24687 53065 24765 53111
rect 24811 53065 24889 53111
rect 24935 53065 25013 53111
rect 25059 53065 25137 53111
rect 25183 53065 25261 53111
rect 25307 53065 25385 53111
rect 25431 53065 25509 53111
rect 25555 53065 25633 53111
rect 25679 53065 25757 53111
rect 25803 53065 25881 53111
rect 25927 53065 26005 53111
rect 26051 53065 26129 53111
rect 26175 53065 26253 53111
rect 26299 53065 26377 53111
rect 26423 53065 26501 53111
rect 26547 53065 26625 53111
rect 26671 53065 26749 53111
rect 26795 53065 26873 53111
rect 26919 53065 26997 53111
rect 27043 53065 27121 53111
rect 27167 53065 27245 53111
rect 27291 53065 27369 53111
rect 27415 53065 27493 53111
rect 27539 53065 27617 53111
rect 27663 53065 27741 53111
rect 27787 53065 27865 53111
rect 27911 53065 27989 53111
rect 28035 53065 28113 53111
rect 28159 53065 28237 53111
rect 28283 53065 28361 53111
rect 28407 53065 28485 53111
rect 28531 53065 28609 53111
rect 28655 53065 28733 53111
rect 28779 53065 28857 53111
rect 28903 53065 28981 53111
rect 29027 53065 29105 53111
rect 29151 53065 29229 53111
rect 29275 53065 29353 53111
rect 29399 53065 29477 53111
rect 29523 53065 29601 53111
rect 29647 53065 29725 53111
rect 29771 53065 29849 53111
rect 29895 53065 29973 53111
rect 30019 53065 30097 53111
rect 30143 53065 30221 53111
rect 30267 53065 30345 53111
rect 30391 53065 30469 53111
rect 30515 53065 30593 53111
rect 30639 53065 30717 53111
rect 30763 53065 30841 53111
rect 30887 53065 30965 53111
rect 31011 53065 31089 53111
rect 31135 53065 31213 53111
rect 31259 53065 31337 53111
rect 31383 53065 31461 53111
rect 31507 53065 31585 53111
rect 31631 53065 31709 53111
rect 31755 53065 31833 53111
rect 31879 53065 31957 53111
rect 32003 53065 32081 53111
rect 32127 53065 32205 53111
rect 32251 53065 32329 53111
rect 32375 53065 32453 53111
rect 32499 53065 32577 53111
rect 32623 53065 32701 53111
rect 32747 53065 32825 53111
rect 32871 53065 32949 53111
rect 32995 53065 33073 53111
rect 33119 53065 33197 53111
rect 33243 53065 33321 53111
rect 33367 53065 33445 53111
rect 33491 53065 33569 53111
rect 33615 53065 33693 53111
rect 33739 53065 33817 53111
rect 33863 53065 33941 53111
rect 33987 53065 34065 53111
rect 34111 53065 34189 53111
rect 34235 53065 34313 53111
rect 34359 53065 34437 53111
rect 34483 53065 34561 53111
rect 34607 53065 34685 53111
rect 34731 53065 34809 53111
rect 34855 53065 34933 53111
rect 34979 53065 35057 53111
rect 35103 53065 35181 53111
rect 35227 53065 35305 53111
rect 35351 53065 35429 53111
rect 35475 53065 35553 53111
rect 35599 53065 35677 53111
rect 35723 53065 35801 53111
rect 35847 53065 35925 53111
rect 35971 53065 36049 53111
rect 36095 53065 36173 53111
rect 36219 53065 36297 53111
rect 36343 53065 36421 53111
rect 36467 53065 36545 53111
rect 36591 53065 36669 53111
rect 36715 53065 36793 53111
rect 36839 53065 36917 53111
rect 36963 53065 37041 53111
rect 37087 53065 37165 53111
rect 37211 53065 37289 53111
rect 37335 53065 37413 53111
rect 37459 53065 37537 53111
rect 37583 53065 37661 53111
rect 37707 53065 37785 53111
rect 37831 53065 37909 53111
rect 37955 53065 38033 53111
rect 38079 53065 38157 53111
rect 38203 53065 38281 53111
rect 38327 53065 38405 53111
rect 38451 53065 38529 53111
rect 38575 53065 38653 53111
rect 38699 53065 38777 53111
rect 38823 53065 38901 53111
rect 38947 53065 39025 53111
rect 39071 53065 39149 53111
rect 39195 53065 39273 53111
rect 39319 53065 39397 53111
rect 39443 53065 39521 53111
rect 39567 53065 39645 53111
rect 39691 53065 39769 53111
rect 39815 53065 39893 53111
rect 39939 53065 40017 53111
rect 40063 53065 40141 53111
rect 40187 53065 40265 53111
rect 40311 53065 40389 53111
rect 40435 53065 40513 53111
rect 40559 53065 40637 53111
rect 40683 53065 40761 53111
rect 40807 53065 40885 53111
rect 40931 53065 41009 53111
rect 41055 53065 41133 53111
rect 41179 53065 41257 53111
rect 41303 53065 41381 53111
rect 41427 53065 41505 53111
rect 41551 53065 41629 53111
rect 41675 53065 41753 53111
rect 41799 53065 41877 53111
rect 41923 53065 42001 53111
rect 42047 53065 42125 53111
rect 42171 53065 42249 53111
rect 42295 53065 42373 53111
rect 42419 53065 42497 53111
rect 42543 53065 42621 53111
rect 42667 53065 42745 53111
rect 42791 53065 42869 53111
rect 42915 53065 42993 53111
rect 43039 53065 43117 53111
rect 43163 53065 43241 53111
rect 43287 53065 43365 53111
rect 43411 53065 43489 53111
rect 43535 53065 43613 53111
rect 43659 53065 43737 53111
rect 43783 53065 43861 53111
rect 43907 53065 43985 53111
rect 44031 53065 44109 53111
rect 44155 53065 44233 53111
rect 44279 53065 44357 53111
rect 44403 53065 44481 53111
rect 44527 53065 44605 53111
rect 44651 53065 44729 53111
rect 44775 53065 44853 53111
rect 44899 53065 44977 53111
rect 45023 53065 45101 53111
rect 45147 53065 45225 53111
rect 45271 53065 45349 53111
rect 45395 53065 45473 53111
rect 45519 53065 45597 53111
rect 45643 53065 45721 53111
rect 45767 53065 45845 53111
rect 45891 53065 45969 53111
rect 46015 53065 46093 53111
rect 46139 53065 46217 53111
rect 46263 53065 46341 53111
rect 46387 53065 46465 53111
rect 46511 53065 46589 53111
rect 46635 53065 46713 53111
rect 46759 53065 46837 53111
rect 46883 53065 46961 53111
rect 47007 53065 47085 53111
rect 47131 53065 47209 53111
rect 47255 53065 47333 53111
rect 47379 53065 47457 53111
rect 47503 53065 47581 53111
rect 47627 53065 47705 53111
rect 47751 53065 47829 53111
rect 47875 53065 47953 53111
rect 47999 53065 48077 53111
rect 48123 53065 48201 53111
rect 48247 53065 48325 53111
rect 48371 53065 48449 53111
rect 48495 53065 48573 53111
rect 48619 53065 48697 53111
rect 48743 53065 48821 53111
rect 48867 53065 48945 53111
rect 48991 53065 49069 53111
rect 49115 53065 49193 53111
rect 49239 53065 49317 53111
rect 49363 53065 49441 53111
rect 49487 53065 49565 53111
rect 49611 53065 49689 53111
rect 49735 53065 49813 53111
rect 49859 53065 49937 53111
rect 49983 53065 50061 53111
rect 50107 53065 50185 53111
rect 50231 53065 50309 53111
rect 50355 53065 50433 53111
rect 50479 53065 50557 53111
rect 50603 53065 50681 53111
rect 50727 53065 50805 53111
rect 50851 53065 50929 53111
rect 50975 53065 51053 53111
rect 51099 53065 51177 53111
rect 51223 53065 51301 53111
rect 51347 53065 51425 53111
rect 51471 53065 51549 53111
rect 51595 53065 51673 53111
rect 51719 53065 51797 53111
rect 51843 53065 51921 53111
rect 51967 53065 52045 53111
rect 52091 53065 52169 53111
rect 52215 53065 52293 53111
rect 52339 53065 52417 53111
rect 52463 53065 52541 53111
rect 52587 53065 52665 53111
rect 52711 53065 52789 53111
rect 52835 53065 52913 53111
rect 52959 53065 53037 53111
rect 53083 53065 53161 53111
rect 53207 53065 53285 53111
rect 53331 53065 53409 53111
rect 53455 53065 53533 53111
rect 53579 53065 53657 53111
rect 53703 53065 53781 53111
rect 53827 53065 53905 53111
rect 53951 53065 54029 53111
rect 54075 53065 54153 53111
rect 54199 53065 54277 53111
rect 54323 53065 54401 53111
rect 54447 53065 54525 53111
rect 54571 53065 54649 53111
rect 54695 53065 54773 53111
rect 54819 53065 54897 53111
rect 54943 53065 55021 53111
rect 55067 53065 55145 53111
rect 55191 53065 55269 53111
rect 55315 53065 55393 53111
rect 55439 53065 55517 53111
rect 55563 53065 55641 53111
rect 55687 53065 55765 53111
rect 55811 53065 55889 53111
rect 55935 53065 56013 53111
rect 56059 53065 56137 53111
rect 56183 53065 56261 53111
rect 56307 53065 56385 53111
rect 56431 53065 56509 53111
rect 56555 53065 56633 53111
rect 56679 53065 56757 53111
rect 56803 53065 56881 53111
rect 56927 53065 57005 53111
rect 57051 53065 57129 53111
rect 57175 53065 57253 53111
rect 57299 53065 57377 53111
rect 57423 53065 57501 53111
rect 57547 53065 57625 53111
rect 57671 53065 57749 53111
rect 57795 53065 57873 53111
rect 57919 53065 57997 53111
rect 58043 53065 58121 53111
rect 58167 53065 58245 53111
rect 58291 53065 58369 53111
rect 58415 53065 58493 53111
rect 58539 53065 58617 53111
rect 58663 53065 58741 53111
rect 58787 53065 58865 53111
rect 58911 53065 58989 53111
rect 59035 53065 59113 53111
rect 59159 53065 59237 53111
rect 59283 53065 59361 53111
rect 59407 53065 59485 53111
rect 59531 53065 59609 53111
rect 59655 53065 59733 53111
rect 59779 53065 59857 53111
rect 59903 53065 59981 53111
rect 60027 53065 60105 53111
rect 60151 53065 60229 53111
rect 60275 53065 60353 53111
rect 60399 53065 60477 53111
rect 60523 53065 60601 53111
rect 60647 53065 60725 53111
rect 60771 53065 60849 53111
rect 60895 53065 60973 53111
rect 61019 53065 61097 53111
rect 61143 53065 61221 53111
rect 61267 53065 61345 53111
rect 61391 53065 61469 53111
rect 61515 53065 61593 53111
rect 61639 53065 61717 53111
rect 61763 53065 61841 53111
rect 61887 53065 61965 53111
rect 62011 53065 62089 53111
rect 62135 53065 62213 53111
rect 62259 53065 62337 53111
rect 62383 53065 62461 53111
rect 62507 53065 62585 53111
rect 62631 53065 62709 53111
rect 62755 53065 62833 53111
rect 62879 53065 62957 53111
rect 63003 53065 63081 53111
rect 63127 53065 63205 53111
rect 63251 53065 63329 53111
rect 63375 53065 63453 53111
rect 63499 53065 63577 53111
rect 63623 53065 63701 53111
rect 63747 53065 63825 53111
rect 63871 53065 63949 53111
rect 63995 53065 64073 53111
rect 64119 53065 64197 53111
rect 64243 53065 64321 53111
rect 64367 53065 64445 53111
rect 64491 53065 64569 53111
rect 64615 53065 64693 53111
rect 64739 53065 64817 53111
rect 64863 53065 64941 53111
rect 64987 53065 65065 53111
rect 65111 53065 65189 53111
rect 65235 53065 65313 53111
rect 65359 53065 65437 53111
rect 65483 53065 65561 53111
rect 65607 53065 65685 53111
rect 65731 53065 65809 53111
rect 65855 53065 65933 53111
rect 65979 53065 66057 53111
rect 66103 53065 66181 53111
rect 66227 53065 66305 53111
rect 66351 53065 66429 53111
rect 66475 53065 66553 53111
rect 66599 53065 66677 53111
rect 66723 53065 66801 53111
rect 66847 53065 66925 53111
rect 66971 53065 67049 53111
rect 67095 53065 67173 53111
rect 67219 53065 67297 53111
rect 67343 53065 67421 53111
rect 67467 53065 67545 53111
rect 67591 53065 67669 53111
rect 67715 53065 67793 53111
rect 67839 53065 67917 53111
rect 67963 53065 68041 53111
rect 68087 53065 68165 53111
rect 68211 53065 68289 53111
rect 68335 53065 68413 53111
rect 68459 53065 68537 53111
rect 68583 53065 68661 53111
rect 68707 53065 68785 53111
rect 68831 53065 68909 53111
rect 68955 53065 69033 53111
rect 69079 53065 69157 53111
rect 69203 53065 69281 53111
rect 69327 53065 69405 53111
rect 69451 53065 69529 53111
rect 69575 53065 69653 53111
rect 69699 53065 69777 53111
rect 69823 53065 69901 53111
rect 69947 53065 70025 53111
rect 70071 53065 70149 53111
rect 70195 53065 70273 53111
rect 70319 53065 70397 53111
rect 70443 53065 70521 53111
rect 70567 53065 70645 53111
rect 70691 53065 70769 53111
rect 70815 53065 70893 53111
rect 70939 53065 71017 53111
rect 71063 53065 71141 53111
rect 71187 53065 71265 53111
rect 71311 53065 71389 53111
rect 71435 53065 71513 53111
rect 71559 53065 71637 53111
rect 71683 53065 71761 53111
rect 71807 53065 71885 53111
rect 71931 53065 72009 53111
rect 72055 53065 72133 53111
rect 72179 53065 72257 53111
rect 72303 53065 72381 53111
rect 72427 53065 72505 53111
rect 72551 53065 72629 53111
rect 72675 53065 72753 53111
rect 72799 53065 72877 53111
rect 72923 53065 73001 53111
rect 73047 53065 73125 53111
rect 73171 53065 73249 53111
rect 73295 53065 73373 53111
rect 73419 53065 73497 53111
rect 73543 53065 73621 53111
rect 73667 53065 73745 53111
rect 73791 53065 73869 53111
rect 73915 53065 73993 53111
rect 74039 53065 74117 53111
rect 74163 53065 74241 53111
rect 74287 53065 74365 53111
rect 74411 53065 74489 53111
rect 74535 53065 74613 53111
rect 74659 53065 74737 53111
rect 74783 53065 74861 53111
rect 74907 53065 74985 53111
rect 75031 53065 75109 53111
rect 75155 53065 75233 53111
rect 75279 53065 75357 53111
rect 75403 53065 75481 53111
rect 75527 53065 75605 53111
rect 75651 53065 75729 53111
rect 75775 53065 75853 53111
rect 75899 53065 75977 53111
rect 76023 53065 76101 53111
rect 76147 53065 76225 53111
rect 76271 53065 76349 53111
rect 76395 53065 76473 53111
rect 76519 53065 76597 53111
rect 76643 53065 76721 53111
rect 76767 53065 76845 53111
rect 76891 53065 76969 53111
rect 77015 53065 77093 53111
rect 77139 53065 77217 53111
rect 77263 53065 77341 53111
rect 77387 53065 77465 53111
rect 77511 53065 77589 53111
rect 77635 53065 77713 53111
rect 77759 53065 77837 53111
rect 77883 53065 77961 53111
rect 78007 53065 78085 53111
rect 78131 53065 78209 53111
rect 78255 53065 78333 53111
rect 78379 53065 78457 53111
rect 78503 53065 78581 53111
rect 78627 53065 78705 53111
rect 78751 53065 78829 53111
rect 78875 53065 78953 53111
rect 78999 53065 79077 53111
rect 79123 53065 79201 53111
rect 79247 53065 79325 53111
rect 79371 53065 79449 53111
rect 79495 53065 79573 53111
rect 79619 53065 79697 53111
rect 79743 53065 79821 53111
rect 79867 53065 79945 53111
rect 79991 53065 80069 53111
rect 80115 53065 80193 53111
rect 80239 53065 80317 53111
rect 80363 53065 80441 53111
rect 80487 53065 80565 53111
rect 80611 53065 80689 53111
rect 80735 53065 80813 53111
rect 80859 53065 80937 53111
rect 80983 53065 81061 53111
rect 81107 53065 81185 53111
rect 81231 53065 81309 53111
rect 81355 53065 81433 53111
rect 81479 53065 81557 53111
rect 81603 53065 81681 53111
rect 81727 53065 81805 53111
rect 81851 53065 81929 53111
rect 81975 53065 82053 53111
rect 82099 53065 82177 53111
rect 82223 53065 82301 53111
rect 82347 53065 82425 53111
rect 82471 53065 82549 53111
rect 82595 53065 82673 53111
rect 82719 53065 82797 53111
rect 82843 53065 82921 53111
rect 82967 53065 83045 53111
rect 83091 53065 83169 53111
rect 83215 53065 83293 53111
rect 83339 53065 83417 53111
rect 83463 53065 83541 53111
rect 83587 53065 83665 53111
rect 83711 53065 83789 53111
rect 83835 53065 83913 53111
rect 83959 53065 84037 53111
rect 84083 53065 84161 53111
rect 84207 53065 84285 53111
rect 84331 53065 84409 53111
rect 84455 53065 84533 53111
rect 84579 53065 84657 53111
rect 84703 53065 84781 53111
rect 84827 53065 84905 53111
rect 84951 53065 85029 53111
rect 85075 53065 85153 53111
rect 85199 53065 85277 53111
rect 85323 53065 85401 53111
rect 85447 53065 85525 53111
rect 85571 53065 85649 53111
rect 85695 53065 85816 53111
rect 70 53046 85816 53065
rect 70 52963 454 53046
rect 70 1117 89 52963
rect 435 1117 454 52963
rect 70 1034 454 1117
rect 85432 52963 85816 53046
rect 85432 1117 85451 52963
rect 85797 1117 85816 52963
rect 85432 1034 85816 1117
rect 70 1015 85816 1034
rect 70 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85816 1015
rect 70 891 85816 969
rect 70 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85816 891
rect 70 767 85816 845
rect 70 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85816 767
rect 70 643 85816 721
rect 70 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85816 643
rect 70 578 85816 597
<< psubdiffcont >>
rect 89 53437 135 53483
rect 213 53437 259 53483
rect 337 53437 383 53483
rect 461 53437 507 53483
rect 585 53437 631 53483
rect 709 53437 755 53483
rect 833 53437 879 53483
rect 957 53437 1003 53483
rect 1081 53437 1127 53483
rect 1205 53437 1251 53483
rect 1329 53437 1375 53483
rect 1453 53437 1499 53483
rect 1577 53437 1623 53483
rect 1701 53437 1747 53483
rect 1825 53437 1871 53483
rect 1949 53437 1995 53483
rect 2073 53437 2119 53483
rect 2197 53437 2243 53483
rect 2321 53437 2367 53483
rect 2445 53437 2491 53483
rect 2569 53437 2615 53483
rect 2693 53437 2739 53483
rect 2817 53437 2863 53483
rect 2941 53437 2987 53483
rect 3065 53437 3111 53483
rect 3189 53437 3235 53483
rect 3313 53437 3359 53483
rect 3437 53437 3483 53483
rect 3561 53437 3607 53483
rect 3685 53437 3731 53483
rect 3809 53437 3855 53483
rect 3933 53437 3979 53483
rect 4057 53437 4103 53483
rect 4181 53437 4227 53483
rect 4305 53437 4351 53483
rect 4429 53437 4475 53483
rect 4553 53437 4599 53483
rect 4677 53437 4723 53483
rect 4801 53437 4847 53483
rect 4925 53437 4971 53483
rect 5049 53437 5095 53483
rect 5173 53437 5219 53483
rect 5297 53437 5343 53483
rect 5421 53437 5467 53483
rect 5545 53437 5591 53483
rect 5669 53437 5715 53483
rect 5793 53437 5839 53483
rect 5917 53437 5963 53483
rect 6041 53437 6087 53483
rect 6165 53437 6211 53483
rect 6289 53437 6335 53483
rect 6413 53437 6459 53483
rect 6537 53437 6583 53483
rect 6661 53437 6707 53483
rect 6785 53437 6831 53483
rect 6909 53437 6955 53483
rect 7033 53437 7079 53483
rect 7157 53437 7203 53483
rect 7281 53437 7327 53483
rect 7405 53437 7451 53483
rect 7529 53437 7575 53483
rect 7653 53437 7699 53483
rect 7777 53437 7823 53483
rect 7901 53437 7947 53483
rect 8025 53437 8071 53483
rect 8149 53437 8195 53483
rect 8273 53437 8319 53483
rect 8397 53437 8443 53483
rect 8521 53437 8567 53483
rect 8645 53437 8691 53483
rect 8769 53437 8815 53483
rect 8893 53437 8939 53483
rect 9017 53437 9063 53483
rect 9141 53437 9187 53483
rect 9265 53437 9311 53483
rect 9389 53437 9435 53483
rect 9513 53437 9559 53483
rect 9637 53437 9683 53483
rect 9761 53437 9807 53483
rect 9885 53437 9931 53483
rect 10009 53437 10055 53483
rect 10133 53437 10179 53483
rect 10257 53437 10303 53483
rect 10381 53437 10427 53483
rect 10505 53437 10551 53483
rect 10629 53437 10675 53483
rect 10753 53437 10799 53483
rect 10877 53437 10923 53483
rect 11001 53437 11047 53483
rect 11125 53437 11171 53483
rect 11249 53437 11295 53483
rect 11373 53437 11419 53483
rect 11497 53437 11543 53483
rect 11621 53437 11667 53483
rect 11745 53437 11791 53483
rect 11869 53437 11915 53483
rect 11993 53437 12039 53483
rect 12117 53437 12163 53483
rect 12241 53437 12287 53483
rect 12365 53437 12411 53483
rect 12489 53437 12535 53483
rect 12613 53437 12659 53483
rect 12737 53437 12783 53483
rect 12861 53437 12907 53483
rect 12985 53437 13031 53483
rect 13109 53437 13155 53483
rect 13233 53437 13279 53483
rect 13357 53437 13403 53483
rect 13481 53437 13527 53483
rect 13605 53437 13651 53483
rect 13729 53437 13775 53483
rect 13853 53437 13899 53483
rect 13977 53437 14023 53483
rect 14101 53437 14147 53483
rect 14225 53437 14271 53483
rect 14349 53437 14395 53483
rect 14473 53437 14519 53483
rect 14597 53437 14643 53483
rect 14721 53437 14767 53483
rect 14845 53437 14891 53483
rect 14969 53437 15015 53483
rect 15093 53437 15139 53483
rect 15217 53437 15263 53483
rect 15341 53437 15387 53483
rect 15465 53437 15511 53483
rect 15589 53437 15635 53483
rect 15713 53437 15759 53483
rect 15837 53437 15883 53483
rect 15961 53437 16007 53483
rect 16085 53437 16131 53483
rect 16209 53437 16255 53483
rect 16333 53437 16379 53483
rect 16457 53437 16503 53483
rect 16581 53437 16627 53483
rect 16705 53437 16751 53483
rect 16829 53437 16875 53483
rect 16953 53437 16999 53483
rect 17077 53437 17123 53483
rect 17201 53437 17247 53483
rect 17325 53437 17371 53483
rect 17449 53437 17495 53483
rect 17573 53437 17619 53483
rect 17697 53437 17743 53483
rect 17821 53437 17867 53483
rect 17945 53437 17991 53483
rect 18069 53437 18115 53483
rect 18193 53437 18239 53483
rect 18317 53437 18363 53483
rect 18441 53437 18487 53483
rect 18565 53437 18611 53483
rect 18689 53437 18735 53483
rect 18813 53437 18859 53483
rect 18937 53437 18983 53483
rect 19061 53437 19107 53483
rect 19185 53437 19231 53483
rect 19309 53437 19355 53483
rect 19433 53437 19479 53483
rect 19557 53437 19603 53483
rect 19681 53437 19727 53483
rect 19805 53437 19851 53483
rect 19929 53437 19975 53483
rect 20053 53437 20099 53483
rect 20177 53437 20223 53483
rect 20301 53437 20347 53483
rect 20425 53437 20471 53483
rect 20549 53437 20595 53483
rect 20673 53437 20719 53483
rect 20797 53437 20843 53483
rect 20921 53437 20967 53483
rect 21045 53437 21091 53483
rect 21169 53437 21215 53483
rect 21293 53437 21339 53483
rect 21417 53437 21463 53483
rect 21541 53437 21587 53483
rect 21665 53437 21711 53483
rect 21789 53437 21835 53483
rect 21913 53437 21959 53483
rect 22037 53437 22083 53483
rect 22161 53437 22207 53483
rect 22285 53437 22331 53483
rect 22409 53437 22455 53483
rect 22533 53437 22579 53483
rect 22657 53437 22703 53483
rect 22781 53437 22827 53483
rect 22905 53437 22951 53483
rect 23029 53437 23075 53483
rect 23153 53437 23199 53483
rect 23277 53437 23323 53483
rect 23401 53437 23447 53483
rect 23525 53437 23571 53483
rect 23649 53437 23695 53483
rect 23773 53437 23819 53483
rect 23897 53437 23943 53483
rect 24021 53437 24067 53483
rect 24145 53437 24191 53483
rect 24269 53437 24315 53483
rect 24393 53437 24439 53483
rect 24517 53437 24563 53483
rect 24641 53437 24687 53483
rect 24765 53437 24811 53483
rect 24889 53437 24935 53483
rect 25013 53437 25059 53483
rect 25137 53437 25183 53483
rect 25261 53437 25307 53483
rect 25385 53437 25431 53483
rect 25509 53437 25555 53483
rect 25633 53437 25679 53483
rect 25757 53437 25803 53483
rect 25881 53437 25927 53483
rect 26005 53437 26051 53483
rect 26129 53437 26175 53483
rect 26253 53437 26299 53483
rect 26377 53437 26423 53483
rect 26501 53437 26547 53483
rect 26625 53437 26671 53483
rect 26749 53437 26795 53483
rect 26873 53437 26919 53483
rect 26997 53437 27043 53483
rect 27121 53437 27167 53483
rect 27245 53437 27291 53483
rect 27369 53437 27415 53483
rect 27493 53437 27539 53483
rect 27617 53437 27663 53483
rect 27741 53437 27787 53483
rect 27865 53437 27911 53483
rect 27989 53437 28035 53483
rect 28113 53437 28159 53483
rect 28237 53437 28283 53483
rect 28361 53437 28407 53483
rect 28485 53437 28531 53483
rect 28609 53437 28655 53483
rect 28733 53437 28779 53483
rect 28857 53437 28903 53483
rect 28981 53437 29027 53483
rect 29105 53437 29151 53483
rect 29229 53437 29275 53483
rect 29353 53437 29399 53483
rect 29477 53437 29523 53483
rect 29601 53437 29647 53483
rect 29725 53437 29771 53483
rect 29849 53437 29895 53483
rect 29973 53437 30019 53483
rect 30097 53437 30143 53483
rect 30221 53437 30267 53483
rect 30345 53437 30391 53483
rect 30469 53437 30515 53483
rect 30593 53437 30639 53483
rect 30717 53437 30763 53483
rect 30841 53437 30887 53483
rect 30965 53437 31011 53483
rect 31089 53437 31135 53483
rect 31213 53437 31259 53483
rect 31337 53437 31383 53483
rect 31461 53437 31507 53483
rect 31585 53437 31631 53483
rect 31709 53437 31755 53483
rect 31833 53437 31879 53483
rect 31957 53437 32003 53483
rect 32081 53437 32127 53483
rect 32205 53437 32251 53483
rect 32329 53437 32375 53483
rect 32453 53437 32499 53483
rect 32577 53437 32623 53483
rect 32701 53437 32747 53483
rect 32825 53437 32871 53483
rect 32949 53437 32995 53483
rect 33073 53437 33119 53483
rect 33197 53437 33243 53483
rect 33321 53437 33367 53483
rect 33445 53437 33491 53483
rect 33569 53437 33615 53483
rect 33693 53437 33739 53483
rect 33817 53437 33863 53483
rect 33941 53437 33987 53483
rect 34065 53437 34111 53483
rect 34189 53437 34235 53483
rect 34313 53437 34359 53483
rect 34437 53437 34483 53483
rect 34561 53437 34607 53483
rect 34685 53437 34731 53483
rect 34809 53437 34855 53483
rect 34933 53437 34979 53483
rect 35057 53437 35103 53483
rect 35181 53437 35227 53483
rect 35305 53437 35351 53483
rect 35429 53437 35475 53483
rect 35553 53437 35599 53483
rect 35677 53437 35723 53483
rect 35801 53437 35847 53483
rect 35925 53437 35971 53483
rect 36049 53437 36095 53483
rect 36173 53437 36219 53483
rect 36297 53437 36343 53483
rect 36421 53437 36467 53483
rect 36545 53437 36591 53483
rect 36669 53437 36715 53483
rect 36793 53437 36839 53483
rect 36917 53437 36963 53483
rect 37041 53437 37087 53483
rect 37165 53437 37211 53483
rect 37289 53437 37335 53483
rect 37413 53437 37459 53483
rect 37537 53437 37583 53483
rect 37661 53437 37707 53483
rect 37785 53437 37831 53483
rect 37909 53437 37955 53483
rect 38033 53437 38079 53483
rect 38157 53437 38203 53483
rect 38281 53437 38327 53483
rect 38405 53437 38451 53483
rect 38529 53437 38575 53483
rect 38653 53437 38699 53483
rect 38777 53437 38823 53483
rect 38901 53437 38947 53483
rect 39025 53437 39071 53483
rect 39149 53437 39195 53483
rect 39273 53437 39319 53483
rect 39397 53437 39443 53483
rect 39521 53437 39567 53483
rect 39645 53437 39691 53483
rect 39769 53437 39815 53483
rect 39893 53437 39939 53483
rect 40017 53437 40063 53483
rect 40141 53437 40187 53483
rect 40265 53437 40311 53483
rect 40389 53437 40435 53483
rect 40513 53437 40559 53483
rect 40637 53437 40683 53483
rect 40761 53437 40807 53483
rect 40885 53437 40931 53483
rect 41009 53437 41055 53483
rect 41133 53437 41179 53483
rect 41257 53437 41303 53483
rect 41381 53437 41427 53483
rect 41505 53437 41551 53483
rect 41629 53437 41675 53483
rect 41753 53437 41799 53483
rect 41877 53437 41923 53483
rect 42001 53437 42047 53483
rect 42125 53437 42171 53483
rect 42249 53437 42295 53483
rect 42373 53437 42419 53483
rect 42497 53437 42543 53483
rect 42621 53437 42667 53483
rect 42745 53437 42791 53483
rect 42869 53437 42915 53483
rect 42993 53437 43039 53483
rect 43117 53437 43163 53483
rect 43241 53437 43287 53483
rect 43365 53437 43411 53483
rect 43489 53437 43535 53483
rect 43613 53437 43659 53483
rect 43737 53437 43783 53483
rect 43861 53437 43907 53483
rect 43985 53437 44031 53483
rect 44109 53437 44155 53483
rect 44233 53437 44279 53483
rect 44357 53437 44403 53483
rect 44481 53437 44527 53483
rect 44605 53437 44651 53483
rect 44729 53437 44775 53483
rect 44853 53437 44899 53483
rect 44977 53437 45023 53483
rect 45101 53437 45147 53483
rect 45225 53437 45271 53483
rect 45349 53437 45395 53483
rect 45473 53437 45519 53483
rect 45597 53437 45643 53483
rect 45721 53437 45767 53483
rect 45845 53437 45891 53483
rect 45969 53437 46015 53483
rect 46093 53437 46139 53483
rect 46217 53437 46263 53483
rect 46341 53437 46387 53483
rect 46465 53437 46511 53483
rect 46589 53437 46635 53483
rect 46713 53437 46759 53483
rect 46837 53437 46883 53483
rect 46961 53437 47007 53483
rect 47085 53437 47131 53483
rect 47209 53437 47255 53483
rect 47333 53437 47379 53483
rect 47457 53437 47503 53483
rect 47581 53437 47627 53483
rect 47705 53437 47751 53483
rect 47829 53437 47875 53483
rect 47953 53437 47999 53483
rect 48077 53437 48123 53483
rect 48201 53437 48247 53483
rect 48325 53437 48371 53483
rect 48449 53437 48495 53483
rect 48573 53437 48619 53483
rect 48697 53437 48743 53483
rect 48821 53437 48867 53483
rect 48945 53437 48991 53483
rect 49069 53437 49115 53483
rect 49193 53437 49239 53483
rect 49317 53437 49363 53483
rect 49441 53437 49487 53483
rect 49565 53437 49611 53483
rect 49689 53437 49735 53483
rect 49813 53437 49859 53483
rect 49937 53437 49983 53483
rect 50061 53437 50107 53483
rect 50185 53437 50231 53483
rect 50309 53437 50355 53483
rect 50433 53437 50479 53483
rect 50557 53437 50603 53483
rect 50681 53437 50727 53483
rect 50805 53437 50851 53483
rect 50929 53437 50975 53483
rect 51053 53437 51099 53483
rect 51177 53437 51223 53483
rect 51301 53437 51347 53483
rect 51425 53437 51471 53483
rect 51549 53437 51595 53483
rect 51673 53437 51719 53483
rect 51797 53437 51843 53483
rect 51921 53437 51967 53483
rect 52045 53437 52091 53483
rect 52169 53437 52215 53483
rect 52293 53437 52339 53483
rect 52417 53437 52463 53483
rect 52541 53437 52587 53483
rect 52665 53437 52711 53483
rect 52789 53437 52835 53483
rect 52913 53437 52959 53483
rect 53037 53437 53083 53483
rect 53161 53437 53207 53483
rect 53285 53437 53331 53483
rect 53409 53437 53455 53483
rect 53533 53437 53579 53483
rect 53657 53437 53703 53483
rect 53781 53437 53827 53483
rect 53905 53437 53951 53483
rect 54029 53437 54075 53483
rect 54153 53437 54199 53483
rect 54277 53437 54323 53483
rect 54401 53437 54447 53483
rect 54525 53437 54571 53483
rect 54649 53437 54695 53483
rect 54773 53437 54819 53483
rect 54897 53437 54943 53483
rect 55021 53437 55067 53483
rect 55145 53437 55191 53483
rect 55269 53437 55315 53483
rect 55393 53437 55439 53483
rect 55517 53437 55563 53483
rect 55641 53437 55687 53483
rect 55765 53437 55811 53483
rect 55889 53437 55935 53483
rect 56013 53437 56059 53483
rect 56137 53437 56183 53483
rect 56261 53437 56307 53483
rect 56385 53437 56431 53483
rect 56509 53437 56555 53483
rect 56633 53437 56679 53483
rect 56757 53437 56803 53483
rect 56881 53437 56927 53483
rect 57005 53437 57051 53483
rect 57129 53437 57175 53483
rect 57253 53437 57299 53483
rect 57377 53437 57423 53483
rect 57501 53437 57547 53483
rect 57625 53437 57671 53483
rect 57749 53437 57795 53483
rect 57873 53437 57919 53483
rect 57997 53437 58043 53483
rect 58121 53437 58167 53483
rect 58245 53437 58291 53483
rect 58369 53437 58415 53483
rect 58493 53437 58539 53483
rect 58617 53437 58663 53483
rect 58741 53437 58787 53483
rect 58865 53437 58911 53483
rect 58989 53437 59035 53483
rect 59113 53437 59159 53483
rect 59237 53437 59283 53483
rect 59361 53437 59407 53483
rect 59485 53437 59531 53483
rect 59609 53437 59655 53483
rect 59733 53437 59779 53483
rect 59857 53437 59903 53483
rect 59981 53437 60027 53483
rect 60105 53437 60151 53483
rect 60229 53437 60275 53483
rect 60353 53437 60399 53483
rect 60477 53437 60523 53483
rect 60601 53437 60647 53483
rect 60725 53437 60771 53483
rect 60849 53437 60895 53483
rect 60973 53437 61019 53483
rect 61097 53437 61143 53483
rect 61221 53437 61267 53483
rect 61345 53437 61391 53483
rect 61469 53437 61515 53483
rect 61593 53437 61639 53483
rect 61717 53437 61763 53483
rect 61841 53437 61887 53483
rect 61965 53437 62011 53483
rect 62089 53437 62135 53483
rect 62213 53437 62259 53483
rect 62337 53437 62383 53483
rect 62461 53437 62507 53483
rect 62585 53437 62631 53483
rect 62709 53437 62755 53483
rect 62833 53437 62879 53483
rect 62957 53437 63003 53483
rect 63081 53437 63127 53483
rect 63205 53437 63251 53483
rect 63329 53437 63375 53483
rect 63453 53437 63499 53483
rect 63577 53437 63623 53483
rect 63701 53437 63747 53483
rect 63825 53437 63871 53483
rect 63949 53437 63995 53483
rect 64073 53437 64119 53483
rect 64197 53437 64243 53483
rect 64321 53437 64367 53483
rect 64445 53437 64491 53483
rect 64569 53437 64615 53483
rect 64693 53437 64739 53483
rect 64817 53437 64863 53483
rect 64941 53437 64987 53483
rect 65065 53437 65111 53483
rect 65189 53437 65235 53483
rect 65313 53437 65359 53483
rect 65437 53437 65483 53483
rect 65561 53437 65607 53483
rect 65685 53437 65731 53483
rect 65809 53437 65855 53483
rect 65933 53437 65979 53483
rect 66057 53437 66103 53483
rect 66181 53437 66227 53483
rect 66305 53437 66351 53483
rect 66429 53437 66475 53483
rect 66553 53437 66599 53483
rect 66677 53437 66723 53483
rect 66801 53437 66847 53483
rect 66925 53437 66971 53483
rect 67049 53437 67095 53483
rect 67173 53437 67219 53483
rect 67297 53437 67343 53483
rect 67421 53437 67467 53483
rect 67545 53437 67591 53483
rect 67669 53437 67715 53483
rect 67793 53437 67839 53483
rect 67917 53437 67963 53483
rect 68041 53437 68087 53483
rect 68165 53437 68211 53483
rect 68289 53437 68335 53483
rect 68413 53437 68459 53483
rect 68537 53437 68583 53483
rect 68661 53437 68707 53483
rect 68785 53437 68831 53483
rect 68909 53437 68955 53483
rect 69033 53437 69079 53483
rect 69157 53437 69203 53483
rect 69281 53437 69327 53483
rect 69405 53437 69451 53483
rect 69529 53437 69575 53483
rect 69653 53437 69699 53483
rect 69777 53437 69823 53483
rect 69901 53437 69947 53483
rect 70025 53437 70071 53483
rect 70149 53437 70195 53483
rect 70273 53437 70319 53483
rect 70397 53437 70443 53483
rect 70521 53437 70567 53483
rect 70645 53437 70691 53483
rect 70769 53437 70815 53483
rect 70893 53437 70939 53483
rect 71017 53437 71063 53483
rect 71141 53437 71187 53483
rect 71265 53437 71311 53483
rect 71389 53437 71435 53483
rect 71513 53437 71559 53483
rect 71637 53437 71683 53483
rect 71761 53437 71807 53483
rect 71885 53437 71931 53483
rect 72009 53437 72055 53483
rect 72133 53437 72179 53483
rect 72257 53437 72303 53483
rect 72381 53437 72427 53483
rect 72505 53437 72551 53483
rect 72629 53437 72675 53483
rect 72753 53437 72799 53483
rect 72877 53437 72923 53483
rect 73001 53437 73047 53483
rect 73125 53437 73171 53483
rect 73249 53437 73295 53483
rect 73373 53437 73419 53483
rect 73497 53437 73543 53483
rect 73621 53437 73667 53483
rect 73745 53437 73791 53483
rect 73869 53437 73915 53483
rect 73993 53437 74039 53483
rect 74117 53437 74163 53483
rect 74241 53437 74287 53483
rect 74365 53437 74411 53483
rect 74489 53437 74535 53483
rect 74613 53437 74659 53483
rect 74737 53437 74783 53483
rect 74861 53437 74907 53483
rect 74985 53437 75031 53483
rect 75109 53437 75155 53483
rect 75233 53437 75279 53483
rect 75357 53437 75403 53483
rect 75481 53437 75527 53483
rect 75605 53437 75651 53483
rect 75729 53437 75775 53483
rect 75853 53437 75899 53483
rect 75977 53437 76023 53483
rect 76101 53437 76147 53483
rect 76225 53437 76271 53483
rect 76349 53437 76395 53483
rect 76473 53437 76519 53483
rect 76597 53437 76643 53483
rect 76721 53437 76767 53483
rect 76845 53437 76891 53483
rect 76969 53437 77015 53483
rect 77093 53437 77139 53483
rect 77217 53437 77263 53483
rect 77341 53437 77387 53483
rect 77465 53437 77511 53483
rect 77589 53437 77635 53483
rect 77713 53437 77759 53483
rect 77837 53437 77883 53483
rect 77961 53437 78007 53483
rect 78085 53437 78131 53483
rect 78209 53437 78255 53483
rect 78333 53437 78379 53483
rect 78457 53437 78503 53483
rect 78581 53437 78627 53483
rect 78705 53437 78751 53483
rect 78829 53437 78875 53483
rect 78953 53437 78999 53483
rect 79077 53437 79123 53483
rect 79201 53437 79247 53483
rect 79325 53437 79371 53483
rect 79449 53437 79495 53483
rect 79573 53437 79619 53483
rect 79697 53437 79743 53483
rect 79821 53437 79867 53483
rect 79945 53437 79991 53483
rect 80069 53437 80115 53483
rect 80193 53437 80239 53483
rect 80317 53437 80363 53483
rect 80441 53437 80487 53483
rect 80565 53437 80611 53483
rect 80689 53437 80735 53483
rect 80813 53437 80859 53483
rect 80937 53437 80983 53483
rect 81061 53437 81107 53483
rect 81185 53437 81231 53483
rect 81309 53437 81355 53483
rect 81433 53437 81479 53483
rect 81557 53437 81603 53483
rect 81681 53437 81727 53483
rect 81805 53437 81851 53483
rect 81929 53437 81975 53483
rect 82053 53437 82099 53483
rect 82177 53437 82223 53483
rect 82301 53437 82347 53483
rect 82425 53437 82471 53483
rect 82549 53437 82595 53483
rect 82673 53437 82719 53483
rect 82797 53437 82843 53483
rect 82921 53437 82967 53483
rect 83045 53437 83091 53483
rect 83169 53437 83215 53483
rect 83293 53437 83339 53483
rect 83417 53437 83463 53483
rect 83541 53437 83587 53483
rect 83665 53437 83711 53483
rect 83789 53437 83835 53483
rect 83913 53437 83959 53483
rect 84037 53437 84083 53483
rect 84161 53437 84207 53483
rect 84285 53437 84331 53483
rect 84409 53437 84455 53483
rect 84533 53437 84579 53483
rect 84657 53437 84703 53483
rect 84781 53437 84827 53483
rect 84905 53437 84951 53483
rect 85029 53437 85075 53483
rect 85153 53437 85199 53483
rect 85277 53437 85323 53483
rect 85401 53437 85447 53483
rect 85525 53437 85571 53483
rect 85649 53437 85695 53483
rect 89 53313 135 53359
rect 213 53313 259 53359
rect 337 53313 383 53359
rect 461 53313 507 53359
rect 585 53313 631 53359
rect 709 53313 755 53359
rect 833 53313 879 53359
rect 957 53313 1003 53359
rect 1081 53313 1127 53359
rect 1205 53313 1251 53359
rect 1329 53313 1375 53359
rect 1453 53313 1499 53359
rect 1577 53313 1623 53359
rect 1701 53313 1747 53359
rect 1825 53313 1871 53359
rect 1949 53313 1995 53359
rect 2073 53313 2119 53359
rect 2197 53313 2243 53359
rect 2321 53313 2367 53359
rect 2445 53313 2491 53359
rect 2569 53313 2615 53359
rect 2693 53313 2739 53359
rect 2817 53313 2863 53359
rect 2941 53313 2987 53359
rect 3065 53313 3111 53359
rect 3189 53313 3235 53359
rect 3313 53313 3359 53359
rect 3437 53313 3483 53359
rect 3561 53313 3607 53359
rect 3685 53313 3731 53359
rect 3809 53313 3855 53359
rect 3933 53313 3979 53359
rect 4057 53313 4103 53359
rect 4181 53313 4227 53359
rect 4305 53313 4351 53359
rect 4429 53313 4475 53359
rect 4553 53313 4599 53359
rect 4677 53313 4723 53359
rect 4801 53313 4847 53359
rect 4925 53313 4971 53359
rect 5049 53313 5095 53359
rect 5173 53313 5219 53359
rect 5297 53313 5343 53359
rect 5421 53313 5467 53359
rect 5545 53313 5591 53359
rect 5669 53313 5715 53359
rect 5793 53313 5839 53359
rect 5917 53313 5963 53359
rect 6041 53313 6087 53359
rect 6165 53313 6211 53359
rect 6289 53313 6335 53359
rect 6413 53313 6459 53359
rect 6537 53313 6583 53359
rect 6661 53313 6707 53359
rect 6785 53313 6831 53359
rect 6909 53313 6955 53359
rect 7033 53313 7079 53359
rect 7157 53313 7203 53359
rect 7281 53313 7327 53359
rect 7405 53313 7451 53359
rect 7529 53313 7575 53359
rect 7653 53313 7699 53359
rect 7777 53313 7823 53359
rect 7901 53313 7947 53359
rect 8025 53313 8071 53359
rect 8149 53313 8195 53359
rect 8273 53313 8319 53359
rect 8397 53313 8443 53359
rect 8521 53313 8567 53359
rect 8645 53313 8691 53359
rect 8769 53313 8815 53359
rect 8893 53313 8939 53359
rect 9017 53313 9063 53359
rect 9141 53313 9187 53359
rect 9265 53313 9311 53359
rect 9389 53313 9435 53359
rect 9513 53313 9559 53359
rect 9637 53313 9683 53359
rect 9761 53313 9807 53359
rect 9885 53313 9931 53359
rect 10009 53313 10055 53359
rect 10133 53313 10179 53359
rect 10257 53313 10303 53359
rect 10381 53313 10427 53359
rect 10505 53313 10551 53359
rect 10629 53313 10675 53359
rect 10753 53313 10799 53359
rect 10877 53313 10923 53359
rect 11001 53313 11047 53359
rect 11125 53313 11171 53359
rect 11249 53313 11295 53359
rect 11373 53313 11419 53359
rect 11497 53313 11543 53359
rect 11621 53313 11667 53359
rect 11745 53313 11791 53359
rect 11869 53313 11915 53359
rect 11993 53313 12039 53359
rect 12117 53313 12163 53359
rect 12241 53313 12287 53359
rect 12365 53313 12411 53359
rect 12489 53313 12535 53359
rect 12613 53313 12659 53359
rect 12737 53313 12783 53359
rect 12861 53313 12907 53359
rect 12985 53313 13031 53359
rect 13109 53313 13155 53359
rect 13233 53313 13279 53359
rect 13357 53313 13403 53359
rect 13481 53313 13527 53359
rect 13605 53313 13651 53359
rect 13729 53313 13775 53359
rect 13853 53313 13899 53359
rect 13977 53313 14023 53359
rect 14101 53313 14147 53359
rect 14225 53313 14271 53359
rect 14349 53313 14395 53359
rect 14473 53313 14519 53359
rect 14597 53313 14643 53359
rect 14721 53313 14767 53359
rect 14845 53313 14891 53359
rect 14969 53313 15015 53359
rect 15093 53313 15139 53359
rect 15217 53313 15263 53359
rect 15341 53313 15387 53359
rect 15465 53313 15511 53359
rect 15589 53313 15635 53359
rect 15713 53313 15759 53359
rect 15837 53313 15883 53359
rect 15961 53313 16007 53359
rect 16085 53313 16131 53359
rect 16209 53313 16255 53359
rect 16333 53313 16379 53359
rect 16457 53313 16503 53359
rect 16581 53313 16627 53359
rect 16705 53313 16751 53359
rect 16829 53313 16875 53359
rect 16953 53313 16999 53359
rect 17077 53313 17123 53359
rect 17201 53313 17247 53359
rect 17325 53313 17371 53359
rect 17449 53313 17495 53359
rect 17573 53313 17619 53359
rect 17697 53313 17743 53359
rect 17821 53313 17867 53359
rect 17945 53313 17991 53359
rect 18069 53313 18115 53359
rect 18193 53313 18239 53359
rect 18317 53313 18363 53359
rect 18441 53313 18487 53359
rect 18565 53313 18611 53359
rect 18689 53313 18735 53359
rect 18813 53313 18859 53359
rect 18937 53313 18983 53359
rect 19061 53313 19107 53359
rect 19185 53313 19231 53359
rect 19309 53313 19355 53359
rect 19433 53313 19479 53359
rect 19557 53313 19603 53359
rect 19681 53313 19727 53359
rect 19805 53313 19851 53359
rect 19929 53313 19975 53359
rect 20053 53313 20099 53359
rect 20177 53313 20223 53359
rect 20301 53313 20347 53359
rect 20425 53313 20471 53359
rect 20549 53313 20595 53359
rect 20673 53313 20719 53359
rect 20797 53313 20843 53359
rect 20921 53313 20967 53359
rect 21045 53313 21091 53359
rect 21169 53313 21215 53359
rect 21293 53313 21339 53359
rect 21417 53313 21463 53359
rect 21541 53313 21587 53359
rect 21665 53313 21711 53359
rect 21789 53313 21835 53359
rect 21913 53313 21959 53359
rect 22037 53313 22083 53359
rect 22161 53313 22207 53359
rect 22285 53313 22331 53359
rect 22409 53313 22455 53359
rect 22533 53313 22579 53359
rect 22657 53313 22703 53359
rect 22781 53313 22827 53359
rect 22905 53313 22951 53359
rect 23029 53313 23075 53359
rect 23153 53313 23199 53359
rect 23277 53313 23323 53359
rect 23401 53313 23447 53359
rect 23525 53313 23571 53359
rect 23649 53313 23695 53359
rect 23773 53313 23819 53359
rect 23897 53313 23943 53359
rect 24021 53313 24067 53359
rect 24145 53313 24191 53359
rect 24269 53313 24315 53359
rect 24393 53313 24439 53359
rect 24517 53313 24563 53359
rect 24641 53313 24687 53359
rect 24765 53313 24811 53359
rect 24889 53313 24935 53359
rect 25013 53313 25059 53359
rect 25137 53313 25183 53359
rect 25261 53313 25307 53359
rect 25385 53313 25431 53359
rect 25509 53313 25555 53359
rect 25633 53313 25679 53359
rect 25757 53313 25803 53359
rect 25881 53313 25927 53359
rect 26005 53313 26051 53359
rect 26129 53313 26175 53359
rect 26253 53313 26299 53359
rect 26377 53313 26423 53359
rect 26501 53313 26547 53359
rect 26625 53313 26671 53359
rect 26749 53313 26795 53359
rect 26873 53313 26919 53359
rect 26997 53313 27043 53359
rect 27121 53313 27167 53359
rect 27245 53313 27291 53359
rect 27369 53313 27415 53359
rect 27493 53313 27539 53359
rect 27617 53313 27663 53359
rect 27741 53313 27787 53359
rect 27865 53313 27911 53359
rect 27989 53313 28035 53359
rect 28113 53313 28159 53359
rect 28237 53313 28283 53359
rect 28361 53313 28407 53359
rect 28485 53313 28531 53359
rect 28609 53313 28655 53359
rect 28733 53313 28779 53359
rect 28857 53313 28903 53359
rect 28981 53313 29027 53359
rect 29105 53313 29151 53359
rect 29229 53313 29275 53359
rect 29353 53313 29399 53359
rect 29477 53313 29523 53359
rect 29601 53313 29647 53359
rect 29725 53313 29771 53359
rect 29849 53313 29895 53359
rect 29973 53313 30019 53359
rect 30097 53313 30143 53359
rect 30221 53313 30267 53359
rect 30345 53313 30391 53359
rect 30469 53313 30515 53359
rect 30593 53313 30639 53359
rect 30717 53313 30763 53359
rect 30841 53313 30887 53359
rect 30965 53313 31011 53359
rect 31089 53313 31135 53359
rect 31213 53313 31259 53359
rect 31337 53313 31383 53359
rect 31461 53313 31507 53359
rect 31585 53313 31631 53359
rect 31709 53313 31755 53359
rect 31833 53313 31879 53359
rect 31957 53313 32003 53359
rect 32081 53313 32127 53359
rect 32205 53313 32251 53359
rect 32329 53313 32375 53359
rect 32453 53313 32499 53359
rect 32577 53313 32623 53359
rect 32701 53313 32747 53359
rect 32825 53313 32871 53359
rect 32949 53313 32995 53359
rect 33073 53313 33119 53359
rect 33197 53313 33243 53359
rect 33321 53313 33367 53359
rect 33445 53313 33491 53359
rect 33569 53313 33615 53359
rect 33693 53313 33739 53359
rect 33817 53313 33863 53359
rect 33941 53313 33987 53359
rect 34065 53313 34111 53359
rect 34189 53313 34235 53359
rect 34313 53313 34359 53359
rect 34437 53313 34483 53359
rect 34561 53313 34607 53359
rect 34685 53313 34731 53359
rect 34809 53313 34855 53359
rect 34933 53313 34979 53359
rect 35057 53313 35103 53359
rect 35181 53313 35227 53359
rect 35305 53313 35351 53359
rect 35429 53313 35475 53359
rect 35553 53313 35599 53359
rect 35677 53313 35723 53359
rect 35801 53313 35847 53359
rect 35925 53313 35971 53359
rect 36049 53313 36095 53359
rect 36173 53313 36219 53359
rect 36297 53313 36343 53359
rect 36421 53313 36467 53359
rect 36545 53313 36591 53359
rect 36669 53313 36715 53359
rect 36793 53313 36839 53359
rect 36917 53313 36963 53359
rect 37041 53313 37087 53359
rect 37165 53313 37211 53359
rect 37289 53313 37335 53359
rect 37413 53313 37459 53359
rect 37537 53313 37583 53359
rect 37661 53313 37707 53359
rect 37785 53313 37831 53359
rect 37909 53313 37955 53359
rect 38033 53313 38079 53359
rect 38157 53313 38203 53359
rect 38281 53313 38327 53359
rect 38405 53313 38451 53359
rect 38529 53313 38575 53359
rect 38653 53313 38699 53359
rect 38777 53313 38823 53359
rect 38901 53313 38947 53359
rect 39025 53313 39071 53359
rect 39149 53313 39195 53359
rect 39273 53313 39319 53359
rect 39397 53313 39443 53359
rect 39521 53313 39567 53359
rect 39645 53313 39691 53359
rect 39769 53313 39815 53359
rect 39893 53313 39939 53359
rect 40017 53313 40063 53359
rect 40141 53313 40187 53359
rect 40265 53313 40311 53359
rect 40389 53313 40435 53359
rect 40513 53313 40559 53359
rect 40637 53313 40683 53359
rect 40761 53313 40807 53359
rect 40885 53313 40931 53359
rect 41009 53313 41055 53359
rect 41133 53313 41179 53359
rect 41257 53313 41303 53359
rect 41381 53313 41427 53359
rect 41505 53313 41551 53359
rect 41629 53313 41675 53359
rect 41753 53313 41799 53359
rect 41877 53313 41923 53359
rect 42001 53313 42047 53359
rect 42125 53313 42171 53359
rect 42249 53313 42295 53359
rect 42373 53313 42419 53359
rect 42497 53313 42543 53359
rect 42621 53313 42667 53359
rect 42745 53313 42791 53359
rect 42869 53313 42915 53359
rect 42993 53313 43039 53359
rect 43117 53313 43163 53359
rect 43241 53313 43287 53359
rect 43365 53313 43411 53359
rect 43489 53313 43535 53359
rect 43613 53313 43659 53359
rect 43737 53313 43783 53359
rect 43861 53313 43907 53359
rect 43985 53313 44031 53359
rect 44109 53313 44155 53359
rect 44233 53313 44279 53359
rect 44357 53313 44403 53359
rect 44481 53313 44527 53359
rect 44605 53313 44651 53359
rect 44729 53313 44775 53359
rect 44853 53313 44899 53359
rect 44977 53313 45023 53359
rect 45101 53313 45147 53359
rect 45225 53313 45271 53359
rect 45349 53313 45395 53359
rect 45473 53313 45519 53359
rect 45597 53313 45643 53359
rect 45721 53313 45767 53359
rect 45845 53313 45891 53359
rect 45969 53313 46015 53359
rect 46093 53313 46139 53359
rect 46217 53313 46263 53359
rect 46341 53313 46387 53359
rect 46465 53313 46511 53359
rect 46589 53313 46635 53359
rect 46713 53313 46759 53359
rect 46837 53313 46883 53359
rect 46961 53313 47007 53359
rect 47085 53313 47131 53359
rect 47209 53313 47255 53359
rect 47333 53313 47379 53359
rect 47457 53313 47503 53359
rect 47581 53313 47627 53359
rect 47705 53313 47751 53359
rect 47829 53313 47875 53359
rect 47953 53313 47999 53359
rect 48077 53313 48123 53359
rect 48201 53313 48247 53359
rect 48325 53313 48371 53359
rect 48449 53313 48495 53359
rect 48573 53313 48619 53359
rect 48697 53313 48743 53359
rect 48821 53313 48867 53359
rect 48945 53313 48991 53359
rect 49069 53313 49115 53359
rect 49193 53313 49239 53359
rect 49317 53313 49363 53359
rect 49441 53313 49487 53359
rect 49565 53313 49611 53359
rect 49689 53313 49735 53359
rect 49813 53313 49859 53359
rect 49937 53313 49983 53359
rect 50061 53313 50107 53359
rect 50185 53313 50231 53359
rect 50309 53313 50355 53359
rect 50433 53313 50479 53359
rect 50557 53313 50603 53359
rect 50681 53313 50727 53359
rect 50805 53313 50851 53359
rect 50929 53313 50975 53359
rect 51053 53313 51099 53359
rect 51177 53313 51223 53359
rect 51301 53313 51347 53359
rect 51425 53313 51471 53359
rect 51549 53313 51595 53359
rect 51673 53313 51719 53359
rect 51797 53313 51843 53359
rect 51921 53313 51967 53359
rect 52045 53313 52091 53359
rect 52169 53313 52215 53359
rect 52293 53313 52339 53359
rect 52417 53313 52463 53359
rect 52541 53313 52587 53359
rect 52665 53313 52711 53359
rect 52789 53313 52835 53359
rect 52913 53313 52959 53359
rect 53037 53313 53083 53359
rect 53161 53313 53207 53359
rect 53285 53313 53331 53359
rect 53409 53313 53455 53359
rect 53533 53313 53579 53359
rect 53657 53313 53703 53359
rect 53781 53313 53827 53359
rect 53905 53313 53951 53359
rect 54029 53313 54075 53359
rect 54153 53313 54199 53359
rect 54277 53313 54323 53359
rect 54401 53313 54447 53359
rect 54525 53313 54571 53359
rect 54649 53313 54695 53359
rect 54773 53313 54819 53359
rect 54897 53313 54943 53359
rect 55021 53313 55067 53359
rect 55145 53313 55191 53359
rect 55269 53313 55315 53359
rect 55393 53313 55439 53359
rect 55517 53313 55563 53359
rect 55641 53313 55687 53359
rect 55765 53313 55811 53359
rect 55889 53313 55935 53359
rect 56013 53313 56059 53359
rect 56137 53313 56183 53359
rect 56261 53313 56307 53359
rect 56385 53313 56431 53359
rect 56509 53313 56555 53359
rect 56633 53313 56679 53359
rect 56757 53313 56803 53359
rect 56881 53313 56927 53359
rect 57005 53313 57051 53359
rect 57129 53313 57175 53359
rect 57253 53313 57299 53359
rect 57377 53313 57423 53359
rect 57501 53313 57547 53359
rect 57625 53313 57671 53359
rect 57749 53313 57795 53359
rect 57873 53313 57919 53359
rect 57997 53313 58043 53359
rect 58121 53313 58167 53359
rect 58245 53313 58291 53359
rect 58369 53313 58415 53359
rect 58493 53313 58539 53359
rect 58617 53313 58663 53359
rect 58741 53313 58787 53359
rect 58865 53313 58911 53359
rect 58989 53313 59035 53359
rect 59113 53313 59159 53359
rect 59237 53313 59283 53359
rect 59361 53313 59407 53359
rect 59485 53313 59531 53359
rect 59609 53313 59655 53359
rect 59733 53313 59779 53359
rect 59857 53313 59903 53359
rect 59981 53313 60027 53359
rect 60105 53313 60151 53359
rect 60229 53313 60275 53359
rect 60353 53313 60399 53359
rect 60477 53313 60523 53359
rect 60601 53313 60647 53359
rect 60725 53313 60771 53359
rect 60849 53313 60895 53359
rect 60973 53313 61019 53359
rect 61097 53313 61143 53359
rect 61221 53313 61267 53359
rect 61345 53313 61391 53359
rect 61469 53313 61515 53359
rect 61593 53313 61639 53359
rect 61717 53313 61763 53359
rect 61841 53313 61887 53359
rect 61965 53313 62011 53359
rect 62089 53313 62135 53359
rect 62213 53313 62259 53359
rect 62337 53313 62383 53359
rect 62461 53313 62507 53359
rect 62585 53313 62631 53359
rect 62709 53313 62755 53359
rect 62833 53313 62879 53359
rect 62957 53313 63003 53359
rect 63081 53313 63127 53359
rect 63205 53313 63251 53359
rect 63329 53313 63375 53359
rect 63453 53313 63499 53359
rect 63577 53313 63623 53359
rect 63701 53313 63747 53359
rect 63825 53313 63871 53359
rect 63949 53313 63995 53359
rect 64073 53313 64119 53359
rect 64197 53313 64243 53359
rect 64321 53313 64367 53359
rect 64445 53313 64491 53359
rect 64569 53313 64615 53359
rect 64693 53313 64739 53359
rect 64817 53313 64863 53359
rect 64941 53313 64987 53359
rect 65065 53313 65111 53359
rect 65189 53313 65235 53359
rect 65313 53313 65359 53359
rect 65437 53313 65483 53359
rect 65561 53313 65607 53359
rect 65685 53313 65731 53359
rect 65809 53313 65855 53359
rect 65933 53313 65979 53359
rect 66057 53313 66103 53359
rect 66181 53313 66227 53359
rect 66305 53313 66351 53359
rect 66429 53313 66475 53359
rect 66553 53313 66599 53359
rect 66677 53313 66723 53359
rect 66801 53313 66847 53359
rect 66925 53313 66971 53359
rect 67049 53313 67095 53359
rect 67173 53313 67219 53359
rect 67297 53313 67343 53359
rect 67421 53313 67467 53359
rect 67545 53313 67591 53359
rect 67669 53313 67715 53359
rect 67793 53313 67839 53359
rect 67917 53313 67963 53359
rect 68041 53313 68087 53359
rect 68165 53313 68211 53359
rect 68289 53313 68335 53359
rect 68413 53313 68459 53359
rect 68537 53313 68583 53359
rect 68661 53313 68707 53359
rect 68785 53313 68831 53359
rect 68909 53313 68955 53359
rect 69033 53313 69079 53359
rect 69157 53313 69203 53359
rect 69281 53313 69327 53359
rect 69405 53313 69451 53359
rect 69529 53313 69575 53359
rect 69653 53313 69699 53359
rect 69777 53313 69823 53359
rect 69901 53313 69947 53359
rect 70025 53313 70071 53359
rect 70149 53313 70195 53359
rect 70273 53313 70319 53359
rect 70397 53313 70443 53359
rect 70521 53313 70567 53359
rect 70645 53313 70691 53359
rect 70769 53313 70815 53359
rect 70893 53313 70939 53359
rect 71017 53313 71063 53359
rect 71141 53313 71187 53359
rect 71265 53313 71311 53359
rect 71389 53313 71435 53359
rect 71513 53313 71559 53359
rect 71637 53313 71683 53359
rect 71761 53313 71807 53359
rect 71885 53313 71931 53359
rect 72009 53313 72055 53359
rect 72133 53313 72179 53359
rect 72257 53313 72303 53359
rect 72381 53313 72427 53359
rect 72505 53313 72551 53359
rect 72629 53313 72675 53359
rect 72753 53313 72799 53359
rect 72877 53313 72923 53359
rect 73001 53313 73047 53359
rect 73125 53313 73171 53359
rect 73249 53313 73295 53359
rect 73373 53313 73419 53359
rect 73497 53313 73543 53359
rect 73621 53313 73667 53359
rect 73745 53313 73791 53359
rect 73869 53313 73915 53359
rect 73993 53313 74039 53359
rect 74117 53313 74163 53359
rect 74241 53313 74287 53359
rect 74365 53313 74411 53359
rect 74489 53313 74535 53359
rect 74613 53313 74659 53359
rect 74737 53313 74783 53359
rect 74861 53313 74907 53359
rect 74985 53313 75031 53359
rect 75109 53313 75155 53359
rect 75233 53313 75279 53359
rect 75357 53313 75403 53359
rect 75481 53313 75527 53359
rect 75605 53313 75651 53359
rect 75729 53313 75775 53359
rect 75853 53313 75899 53359
rect 75977 53313 76023 53359
rect 76101 53313 76147 53359
rect 76225 53313 76271 53359
rect 76349 53313 76395 53359
rect 76473 53313 76519 53359
rect 76597 53313 76643 53359
rect 76721 53313 76767 53359
rect 76845 53313 76891 53359
rect 76969 53313 77015 53359
rect 77093 53313 77139 53359
rect 77217 53313 77263 53359
rect 77341 53313 77387 53359
rect 77465 53313 77511 53359
rect 77589 53313 77635 53359
rect 77713 53313 77759 53359
rect 77837 53313 77883 53359
rect 77961 53313 78007 53359
rect 78085 53313 78131 53359
rect 78209 53313 78255 53359
rect 78333 53313 78379 53359
rect 78457 53313 78503 53359
rect 78581 53313 78627 53359
rect 78705 53313 78751 53359
rect 78829 53313 78875 53359
rect 78953 53313 78999 53359
rect 79077 53313 79123 53359
rect 79201 53313 79247 53359
rect 79325 53313 79371 53359
rect 79449 53313 79495 53359
rect 79573 53313 79619 53359
rect 79697 53313 79743 53359
rect 79821 53313 79867 53359
rect 79945 53313 79991 53359
rect 80069 53313 80115 53359
rect 80193 53313 80239 53359
rect 80317 53313 80363 53359
rect 80441 53313 80487 53359
rect 80565 53313 80611 53359
rect 80689 53313 80735 53359
rect 80813 53313 80859 53359
rect 80937 53313 80983 53359
rect 81061 53313 81107 53359
rect 81185 53313 81231 53359
rect 81309 53313 81355 53359
rect 81433 53313 81479 53359
rect 81557 53313 81603 53359
rect 81681 53313 81727 53359
rect 81805 53313 81851 53359
rect 81929 53313 81975 53359
rect 82053 53313 82099 53359
rect 82177 53313 82223 53359
rect 82301 53313 82347 53359
rect 82425 53313 82471 53359
rect 82549 53313 82595 53359
rect 82673 53313 82719 53359
rect 82797 53313 82843 53359
rect 82921 53313 82967 53359
rect 83045 53313 83091 53359
rect 83169 53313 83215 53359
rect 83293 53313 83339 53359
rect 83417 53313 83463 53359
rect 83541 53313 83587 53359
rect 83665 53313 83711 53359
rect 83789 53313 83835 53359
rect 83913 53313 83959 53359
rect 84037 53313 84083 53359
rect 84161 53313 84207 53359
rect 84285 53313 84331 53359
rect 84409 53313 84455 53359
rect 84533 53313 84579 53359
rect 84657 53313 84703 53359
rect 84781 53313 84827 53359
rect 84905 53313 84951 53359
rect 85029 53313 85075 53359
rect 85153 53313 85199 53359
rect 85277 53313 85323 53359
rect 85401 53313 85447 53359
rect 85525 53313 85571 53359
rect 85649 53313 85695 53359
rect 89 53189 135 53235
rect 213 53189 259 53235
rect 337 53189 383 53235
rect 461 53189 507 53235
rect 585 53189 631 53235
rect 709 53189 755 53235
rect 833 53189 879 53235
rect 957 53189 1003 53235
rect 1081 53189 1127 53235
rect 1205 53189 1251 53235
rect 1329 53189 1375 53235
rect 1453 53189 1499 53235
rect 1577 53189 1623 53235
rect 1701 53189 1747 53235
rect 1825 53189 1871 53235
rect 1949 53189 1995 53235
rect 2073 53189 2119 53235
rect 2197 53189 2243 53235
rect 2321 53189 2367 53235
rect 2445 53189 2491 53235
rect 2569 53189 2615 53235
rect 2693 53189 2739 53235
rect 2817 53189 2863 53235
rect 2941 53189 2987 53235
rect 3065 53189 3111 53235
rect 3189 53189 3235 53235
rect 3313 53189 3359 53235
rect 3437 53189 3483 53235
rect 3561 53189 3607 53235
rect 3685 53189 3731 53235
rect 3809 53189 3855 53235
rect 3933 53189 3979 53235
rect 4057 53189 4103 53235
rect 4181 53189 4227 53235
rect 4305 53189 4351 53235
rect 4429 53189 4475 53235
rect 4553 53189 4599 53235
rect 4677 53189 4723 53235
rect 4801 53189 4847 53235
rect 4925 53189 4971 53235
rect 5049 53189 5095 53235
rect 5173 53189 5219 53235
rect 5297 53189 5343 53235
rect 5421 53189 5467 53235
rect 5545 53189 5591 53235
rect 5669 53189 5715 53235
rect 5793 53189 5839 53235
rect 5917 53189 5963 53235
rect 6041 53189 6087 53235
rect 6165 53189 6211 53235
rect 6289 53189 6335 53235
rect 6413 53189 6459 53235
rect 6537 53189 6583 53235
rect 6661 53189 6707 53235
rect 6785 53189 6831 53235
rect 6909 53189 6955 53235
rect 7033 53189 7079 53235
rect 7157 53189 7203 53235
rect 7281 53189 7327 53235
rect 7405 53189 7451 53235
rect 7529 53189 7575 53235
rect 7653 53189 7699 53235
rect 7777 53189 7823 53235
rect 7901 53189 7947 53235
rect 8025 53189 8071 53235
rect 8149 53189 8195 53235
rect 8273 53189 8319 53235
rect 8397 53189 8443 53235
rect 8521 53189 8567 53235
rect 8645 53189 8691 53235
rect 8769 53189 8815 53235
rect 8893 53189 8939 53235
rect 9017 53189 9063 53235
rect 9141 53189 9187 53235
rect 9265 53189 9311 53235
rect 9389 53189 9435 53235
rect 9513 53189 9559 53235
rect 9637 53189 9683 53235
rect 9761 53189 9807 53235
rect 9885 53189 9931 53235
rect 10009 53189 10055 53235
rect 10133 53189 10179 53235
rect 10257 53189 10303 53235
rect 10381 53189 10427 53235
rect 10505 53189 10551 53235
rect 10629 53189 10675 53235
rect 10753 53189 10799 53235
rect 10877 53189 10923 53235
rect 11001 53189 11047 53235
rect 11125 53189 11171 53235
rect 11249 53189 11295 53235
rect 11373 53189 11419 53235
rect 11497 53189 11543 53235
rect 11621 53189 11667 53235
rect 11745 53189 11791 53235
rect 11869 53189 11915 53235
rect 11993 53189 12039 53235
rect 12117 53189 12163 53235
rect 12241 53189 12287 53235
rect 12365 53189 12411 53235
rect 12489 53189 12535 53235
rect 12613 53189 12659 53235
rect 12737 53189 12783 53235
rect 12861 53189 12907 53235
rect 12985 53189 13031 53235
rect 13109 53189 13155 53235
rect 13233 53189 13279 53235
rect 13357 53189 13403 53235
rect 13481 53189 13527 53235
rect 13605 53189 13651 53235
rect 13729 53189 13775 53235
rect 13853 53189 13899 53235
rect 13977 53189 14023 53235
rect 14101 53189 14147 53235
rect 14225 53189 14271 53235
rect 14349 53189 14395 53235
rect 14473 53189 14519 53235
rect 14597 53189 14643 53235
rect 14721 53189 14767 53235
rect 14845 53189 14891 53235
rect 14969 53189 15015 53235
rect 15093 53189 15139 53235
rect 15217 53189 15263 53235
rect 15341 53189 15387 53235
rect 15465 53189 15511 53235
rect 15589 53189 15635 53235
rect 15713 53189 15759 53235
rect 15837 53189 15883 53235
rect 15961 53189 16007 53235
rect 16085 53189 16131 53235
rect 16209 53189 16255 53235
rect 16333 53189 16379 53235
rect 16457 53189 16503 53235
rect 16581 53189 16627 53235
rect 16705 53189 16751 53235
rect 16829 53189 16875 53235
rect 16953 53189 16999 53235
rect 17077 53189 17123 53235
rect 17201 53189 17247 53235
rect 17325 53189 17371 53235
rect 17449 53189 17495 53235
rect 17573 53189 17619 53235
rect 17697 53189 17743 53235
rect 17821 53189 17867 53235
rect 17945 53189 17991 53235
rect 18069 53189 18115 53235
rect 18193 53189 18239 53235
rect 18317 53189 18363 53235
rect 18441 53189 18487 53235
rect 18565 53189 18611 53235
rect 18689 53189 18735 53235
rect 18813 53189 18859 53235
rect 18937 53189 18983 53235
rect 19061 53189 19107 53235
rect 19185 53189 19231 53235
rect 19309 53189 19355 53235
rect 19433 53189 19479 53235
rect 19557 53189 19603 53235
rect 19681 53189 19727 53235
rect 19805 53189 19851 53235
rect 19929 53189 19975 53235
rect 20053 53189 20099 53235
rect 20177 53189 20223 53235
rect 20301 53189 20347 53235
rect 20425 53189 20471 53235
rect 20549 53189 20595 53235
rect 20673 53189 20719 53235
rect 20797 53189 20843 53235
rect 20921 53189 20967 53235
rect 21045 53189 21091 53235
rect 21169 53189 21215 53235
rect 21293 53189 21339 53235
rect 21417 53189 21463 53235
rect 21541 53189 21587 53235
rect 21665 53189 21711 53235
rect 21789 53189 21835 53235
rect 21913 53189 21959 53235
rect 22037 53189 22083 53235
rect 22161 53189 22207 53235
rect 22285 53189 22331 53235
rect 22409 53189 22455 53235
rect 22533 53189 22579 53235
rect 22657 53189 22703 53235
rect 22781 53189 22827 53235
rect 22905 53189 22951 53235
rect 23029 53189 23075 53235
rect 23153 53189 23199 53235
rect 23277 53189 23323 53235
rect 23401 53189 23447 53235
rect 23525 53189 23571 53235
rect 23649 53189 23695 53235
rect 23773 53189 23819 53235
rect 23897 53189 23943 53235
rect 24021 53189 24067 53235
rect 24145 53189 24191 53235
rect 24269 53189 24315 53235
rect 24393 53189 24439 53235
rect 24517 53189 24563 53235
rect 24641 53189 24687 53235
rect 24765 53189 24811 53235
rect 24889 53189 24935 53235
rect 25013 53189 25059 53235
rect 25137 53189 25183 53235
rect 25261 53189 25307 53235
rect 25385 53189 25431 53235
rect 25509 53189 25555 53235
rect 25633 53189 25679 53235
rect 25757 53189 25803 53235
rect 25881 53189 25927 53235
rect 26005 53189 26051 53235
rect 26129 53189 26175 53235
rect 26253 53189 26299 53235
rect 26377 53189 26423 53235
rect 26501 53189 26547 53235
rect 26625 53189 26671 53235
rect 26749 53189 26795 53235
rect 26873 53189 26919 53235
rect 26997 53189 27043 53235
rect 27121 53189 27167 53235
rect 27245 53189 27291 53235
rect 27369 53189 27415 53235
rect 27493 53189 27539 53235
rect 27617 53189 27663 53235
rect 27741 53189 27787 53235
rect 27865 53189 27911 53235
rect 27989 53189 28035 53235
rect 28113 53189 28159 53235
rect 28237 53189 28283 53235
rect 28361 53189 28407 53235
rect 28485 53189 28531 53235
rect 28609 53189 28655 53235
rect 28733 53189 28779 53235
rect 28857 53189 28903 53235
rect 28981 53189 29027 53235
rect 29105 53189 29151 53235
rect 29229 53189 29275 53235
rect 29353 53189 29399 53235
rect 29477 53189 29523 53235
rect 29601 53189 29647 53235
rect 29725 53189 29771 53235
rect 29849 53189 29895 53235
rect 29973 53189 30019 53235
rect 30097 53189 30143 53235
rect 30221 53189 30267 53235
rect 30345 53189 30391 53235
rect 30469 53189 30515 53235
rect 30593 53189 30639 53235
rect 30717 53189 30763 53235
rect 30841 53189 30887 53235
rect 30965 53189 31011 53235
rect 31089 53189 31135 53235
rect 31213 53189 31259 53235
rect 31337 53189 31383 53235
rect 31461 53189 31507 53235
rect 31585 53189 31631 53235
rect 31709 53189 31755 53235
rect 31833 53189 31879 53235
rect 31957 53189 32003 53235
rect 32081 53189 32127 53235
rect 32205 53189 32251 53235
rect 32329 53189 32375 53235
rect 32453 53189 32499 53235
rect 32577 53189 32623 53235
rect 32701 53189 32747 53235
rect 32825 53189 32871 53235
rect 32949 53189 32995 53235
rect 33073 53189 33119 53235
rect 33197 53189 33243 53235
rect 33321 53189 33367 53235
rect 33445 53189 33491 53235
rect 33569 53189 33615 53235
rect 33693 53189 33739 53235
rect 33817 53189 33863 53235
rect 33941 53189 33987 53235
rect 34065 53189 34111 53235
rect 34189 53189 34235 53235
rect 34313 53189 34359 53235
rect 34437 53189 34483 53235
rect 34561 53189 34607 53235
rect 34685 53189 34731 53235
rect 34809 53189 34855 53235
rect 34933 53189 34979 53235
rect 35057 53189 35103 53235
rect 35181 53189 35227 53235
rect 35305 53189 35351 53235
rect 35429 53189 35475 53235
rect 35553 53189 35599 53235
rect 35677 53189 35723 53235
rect 35801 53189 35847 53235
rect 35925 53189 35971 53235
rect 36049 53189 36095 53235
rect 36173 53189 36219 53235
rect 36297 53189 36343 53235
rect 36421 53189 36467 53235
rect 36545 53189 36591 53235
rect 36669 53189 36715 53235
rect 36793 53189 36839 53235
rect 36917 53189 36963 53235
rect 37041 53189 37087 53235
rect 37165 53189 37211 53235
rect 37289 53189 37335 53235
rect 37413 53189 37459 53235
rect 37537 53189 37583 53235
rect 37661 53189 37707 53235
rect 37785 53189 37831 53235
rect 37909 53189 37955 53235
rect 38033 53189 38079 53235
rect 38157 53189 38203 53235
rect 38281 53189 38327 53235
rect 38405 53189 38451 53235
rect 38529 53189 38575 53235
rect 38653 53189 38699 53235
rect 38777 53189 38823 53235
rect 38901 53189 38947 53235
rect 39025 53189 39071 53235
rect 39149 53189 39195 53235
rect 39273 53189 39319 53235
rect 39397 53189 39443 53235
rect 39521 53189 39567 53235
rect 39645 53189 39691 53235
rect 39769 53189 39815 53235
rect 39893 53189 39939 53235
rect 40017 53189 40063 53235
rect 40141 53189 40187 53235
rect 40265 53189 40311 53235
rect 40389 53189 40435 53235
rect 40513 53189 40559 53235
rect 40637 53189 40683 53235
rect 40761 53189 40807 53235
rect 40885 53189 40931 53235
rect 41009 53189 41055 53235
rect 41133 53189 41179 53235
rect 41257 53189 41303 53235
rect 41381 53189 41427 53235
rect 41505 53189 41551 53235
rect 41629 53189 41675 53235
rect 41753 53189 41799 53235
rect 41877 53189 41923 53235
rect 42001 53189 42047 53235
rect 42125 53189 42171 53235
rect 42249 53189 42295 53235
rect 42373 53189 42419 53235
rect 42497 53189 42543 53235
rect 42621 53189 42667 53235
rect 42745 53189 42791 53235
rect 42869 53189 42915 53235
rect 42993 53189 43039 53235
rect 43117 53189 43163 53235
rect 43241 53189 43287 53235
rect 43365 53189 43411 53235
rect 43489 53189 43535 53235
rect 43613 53189 43659 53235
rect 43737 53189 43783 53235
rect 43861 53189 43907 53235
rect 43985 53189 44031 53235
rect 44109 53189 44155 53235
rect 44233 53189 44279 53235
rect 44357 53189 44403 53235
rect 44481 53189 44527 53235
rect 44605 53189 44651 53235
rect 44729 53189 44775 53235
rect 44853 53189 44899 53235
rect 44977 53189 45023 53235
rect 45101 53189 45147 53235
rect 45225 53189 45271 53235
rect 45349 53189 45395 53235
rect 45473 53189 45519 53235
rect 45597 53189 45643 53235
rect 45721 53189 45767 53235
rect 45845 53189 45891 53235
rect 45969 53189 46015 53235
rect 46093 53189 46139 53235
rect 46217 53189 46263 53235
rect 46341 53189 46387 53235
rect 46465 53189 46511 53235
rect 46589 53189 46635 53235
rect 46713 53189 46759 53235
rect 46837 53189 46883 53235
rect 46961 53189 47007 53235
rect 47085 53189 47131 53235
rect 47209 53189 47255 53235
rect 47333 53189 47379 53235
rect 47457 53189 47503 53235
rect 47581 53189 47627 53235
rect 47705 53189 47751 53235
rect 47829 53189 47875 53235
rect 47953 53189 47999 53235
rect 48077 53189 48123 53235
rect 48201 53189 48247 53235
rect 48325 53189 48371 53235
rect 48449 53189 48495 53235
rect 48573 53189 48619 53235
rect 48697 53189 48743 53235
rect 48821 53189 48867 53235
rect 48945 53189 48991 53235
rect 49069 53189 49115 53235
rect 49193 53189 49239 53235
rect 49317 53189 49363 53235
rect 49441 53189 49487 53235
rect 49565 53189 49611 53235
rect 49689 53189 49735 53235
rect 49813 53189 49859 53235
rect 49937 53189 49983 53235
rect 50061 53189 50107 53235
rect 50185 53189 50231 53235
rect 50309 53189 50355 53235
rect 50433 53189 50479 53235
rect 50557 53189 50603 53235
rect 50681 53189 50727 53235
rect 50805 53189 50851 53235
rect 50929 53189 50975 53235
rect 51053 53189 51099 53235
rect 51177 53189 51223 53235
rect 51301 53189 51347 53235
rect 51425 53189 51471 53235
rect 51549 53189 51595 53235
rect 51673 53189 51719 53235
rect 51797 53189 51843 53235
rect 51921 53189 51967 53235
rect 52045 53189 52091 53235
rect 52169 53189 52215 53235
rect 52293 53189 52339 53235
rect 52417 53189 52463 53235
rect 52541 53189 52587 53235
rect 52665 53189 52711 53235
rect 52789 53189 52835 53235
rect 52913 53189 52959 53235
rect 53037 53189 53083 53235
rect 53161 53189 53207 53235
rect 53285 53189 53331 53235
rect 53409 53189 53455 53235
rect 53533 53189 53579 53235
rect 53657 53189 53703 53235
rect 53781 53189 53827 53235
rect 53905 53189 53951 53235
rect 54029 53189 54075 53235
rect 54153 53189 54199 53235
rect 54277 53189 54323 53235
rect 54401 53189 54447 53235
rect 54525 53189 54571 53235
rect 54649 53189 54695 53235
rect 54773 53189 54819 53235
rect 54897 53189 54943 53235
rect 55021 53189 55067 53235
rect 55145 53189 55191 53235
rect 55269 53189 55315 53235
rect 55393 53189 55439 53235
rect 55517 53189 55563 53235
rect 55641 53189 55687 53235
rect 55765 53189 55811 53235
rect 55889 53189 55935 53235
rect 56013 53189 56059 53235
rect 56137 53189 56183 53235
rect 56261 53189 56307 53235
rect 56385 53189 56431 53235
rect 56509 53189 56555 53235
rect 56633 53189 56679 53235
rect 56757 53189 56803 53235
rect 56881 53189 56927 53235
rect 57005 53189 57051 53235
rect 57129 53189 57175 53235
rect 57253 53189 57299 53235
rect 57377 53189 57423 53235
rect 57501 53189 57547 53235
rect 57625 53189 57671 53235
rect 57749 53189 57795 53235
rect 57873 53189 57919 53235
rect 57997 53189 58043 53235
rect 58121 53189 58167 53235
rect 58245 53189 58291 53235
rect 58369 53189 58415 53235
rect 58493 53189 58539 53235
rect 58617 53189 58663 53235
rect 58741 53189 58787 53235
rect 58865 53189 58911 53235
rect 58989 53189 59035 53235
rect 59113 53189 59159 53235
rect 59237 53189 59283 53235
rect 59361 53189 59407 53235
rect 59485 53189 59531 53235
rect 59609 53189 59655 53235
rect 59733 53189 59779 53235
rect 59857 53189 59903 53235
rect 59981 53189 60027 53235
rect 60105 53189 60151 53235
rect 60229 53189 60275 53235
rect 60353 53189 60399 53235
rect 60477 53189 60523 53235
rect 60601 53189 60647 53235
rect 60725 53189 60771 53235
rect 60849 53189 60895 53235
rect 60973 53189 61019 53235
rect 61097 53189 61143 53235
rect 61221 53189 61267 53235
rect 61345 53189 61391 53235
rect 61469 53189 61515 53235
rect 61593 53189 61639 53235
rect 61717 53189 61763 53235
rect 61841 53189 61887 53235
rect 61965 53189 62011 53235
rect 62089 53189 62135 53235
rect 62213 53189 62259 53235
rect 62337 53189 62383 53235
rect 62461 53189 62507 53235
rect 62585 53189 62631 53235
rect 62709 53189 62755 53235
rect 62833 53189 62879 53235
rect 62957 53189 63003 53235
rect 63081 53189 63127 53235
rect 63205 53189 63251 53235
rect 63329 53189 63375 53235
rect 63453 53189 63499 53235
rect 63577 53189 63623 53235
rect 63701 53189 63747 53235
rect 63825 53189 63871 53235
rect 63949 53189 63995 53235
rect 64073 53189 64119 53235
rect 64197 53189 64243 53235
rect 64321 53189 64367 53235
rect 64445 53189 64491 53235
rect 64569 53189 64615 53235
rect 64693 53189 64739 53235
rect 64817 53189 64863 53235
rect 64941 53189 64987 53235
rect 65065 53189 65111 53235
rect 65189 53189 65235 53235
rect 65313 53189 65359 53235
rect 65437 53189 65483 53235
rect 65561 53189 65607 53235
rect 65685 53189 65731 53235
rect 65809 53189 65855 53235
rect 65933 53189 65979 53235
rect 66057 53189 66103 53235
rect 66181 53189 66227 53235
rect 66305 53189 66351 53235
rect 66429 53189 66475 53235
rect 66553 53189 66599 53235
rect 66677 53189 66723 53235
rect 66801 53189 66847 53235
rect 66925 53189 66971 53235
rect 67049 53189 67095 53235
rect 67173 53189 67219 53235
rect 67297 53189 67343 53235
rect 67421 53189 67467 53235
rect 67545 53189 67591 53235
rect 67669 53189 67715 53235
rect 67793 53189 67839 53235
rect 67917 53189 67963 53235
rect 68041 53189 68087 53235
rect 68165 53189 68211 53235
rect 68289 53189 68335 53235
rect 68413 53189 68459 53235
rect 68537 53189 68583 53235
rect 68661 53189 68707 53235
rect 68785 53189 68831 53235
rect 68909 53189 68955 53235
rect 69033 53189 69079 53235
rect 69157 53189 69203 53235
rect 69281 53189 69327 53235
rect 69405 53189 69451 53235
rect 69529 53189 69575 53235
rect 69653 53189 69699 53235
rect 69777 53189 69823 53235
rect 69901 53189 69947 53235
rect 70025 53189 70071 53235
rect 70149 53189 70195 53235
rect 70273 53189 70319 53235
rect 70397 53189 70443 53235
rect 70521 53189 70567 53235
rect 70645 53189 70691 53235
rect 70769 53189 70815 53235
rect 70893 53189 70939 53235
rect 71017 53189 71063 53235
rect 71141 53189 71187 53235
rect 71265 53189 71311 53235
rect 71389 53189 71435 53235
rect 71513 53189 71559 53235
rect 71637 53189 71683 53235
rect 71761 53189 71807 53235
rect 71885 53189 71931 53235
rect 72009 53189 72055 53235
rect 72133 53189 72179 53235
rect 72257 53189 72303 53235
rect 72381 53189 72427 53235
rect 72505 53189 72551 53235
rect 72629 53189 72675 53235
rect 72753 53189 72799 53235
rect 72877 53189 72923 53235
rect 73001 53189 73047 53235
rect 73125 53189 73171 53235
rect 73249 53189 73295 53235
rect 73373 53189 73419 53235
rect 73497 53189 73543 53235
rect 73621 53189 73667 53235
rect 73745 53189 73791 53235
rect 73869 53189 73915 53235
rect 73993 53189 74039 53235
rect 74117 53189 74163 53235
rect 74241 53189 74287 53235
rect 74365 53189 74411 53235
rect 74489 53189 74535 53235
rect 74613 53189 74659 53235
rect 74737 53189 74783 53235
rect 74861 53189 74907 53235
rect 74985 53189 75031 53235
rect 75109 53189 75155 53235
rect 75233 53189 75279 53235
rect 75357 53189 75403 53235
rect 75481 53189 75527 53235
rect 75605 53189 75651 53235
rect 75729 53189 75775 53235
rect 75853 53189 75899 53235
rect 75977 53189 76023 53235
rect 76101 53189 76147 53235
rect 76225 53189 76271 53235
rect 76349 53189 76395 53235
rect 76473 53189 76519 53235
rect 76597 53189 76643 53235
rect 76721 53189 76767 53235
rect 76845 53189 76891 53235
rect 76969 53189 77015 53235
rect 77093 53189 77139 53235
rect 77217 53189 77263 53235
rect 77341 53189 77387 53235
rect 77465 53189 77511 53235
rect 77589 53189 77635 53235
rect 77713 53189 77759 53235
rect 77837 53189 77883 53235
rect 77961 53189 78007 53235
rect 78085 53189 78131 53235
rect 78209 53189 78255 53235
rect 78333 53189 78379 53235
rect 78457 53189 78503 53235
rect 78581 53189 78627 53235
rect 78705 53189 78751 53235
rect 78829 53189 78875 53235
rect 78953 53189 78999 53235
rect 79077 53189 79123 53235
rect 79201 53189 79247 53235
rect 79325 53189 79371 53235
rect 79449 53189 79495 53235
rect 79573 53189 79619 53235
rect 79697 53189 79743 53235
rect 79821 53189 79867 53235
rect 79945 53189 79991 53235
rect 80069 53189 80115 53235
rect 80193 53189 80239 53235
rect 80317 53189 80363 53235
rect 80441 53189 80487 53235
rect 80565 53189 80611 53235
rect 80689 53189 80735 53235
rect 80813 53189 80859 53235
rect 80937 53189 80983 53235
rect 81061 53189 81107 53235
rect 81185 53189 81231 53235
rect 81309 53189 81355 53235
rect 81433 53189 81479 53235
rect 81557 53189 81603 53235
rect 81681 53189 81727 53235
rect 81805 53189 81851 53235
rect 81929 53189 81975 53235
rect 82053 53189 82099 53235
rect 82177 53189 82223 53235
rect 82301 53189 82347 53235
rect 82425 53189 82471 53235
rect 82549 53189 82595 53235
rect 82673 53189 82719 53235
rect 82797 53189 82843 53235
rect 82921 53189 82967 53235
rect 83045 53189 83091 53235
rect 83169 53189 83215 53235
rect 83293 53189 83339 53235
rect 83417 53189 83463 53235
rect 83541 53189 83587 53235
rect 83665 53189 83711 53235
rect 83789 53189 83835 53235
rect 83913 53189 83959 53235
rect 84037 53189 84083 53235
rect 84161 53189 84207 53235
rect 84285 53189 84331 53235
rect 84409 53189 84455 53235
rect 84533 53189 84579 53235
rect 84657 53189 84703 53235
rect 84781 53189 84827 53235
rect 84905 53189 84951 53235
rect 85029 53189 85075 53235
rect 85153 53189 85199 53235
rect 85277 53189 85323 53235
rect 85401 53189 85447 53235
rect 85525 53189 85571 53235
rect 85649 53189 85695 53235
rect 89 53065 135 53111
rect 213 53065 259 53111
rect 337 53065 383 53111
rect 461 53065 507 53111
rect 585 53065 631 53111
rect 709 53065 755 53111
rect 833 53065 879 53111
rect 957 53065 1003 53111
rect 1081 53065 1127 53111
rect 1205 53065 1251 53111
rect 1329 53065 1375 53111
rect 1453 53065 1499 53111
rect 1577 53065 1623 53111
rect 1701 53065 1747 53111
rect 1825 53065 1871 53111
rect 1949 53065 1995 53111
rect 2073 53065 2119 53111
rect 2197 53065 2243 53111
rect 2321 53065 2367 53111
rect 2445 53065 2491 53111
rect 2569 53065 2615 53111
rect 2693 53065 2739 53111
rect 2817 53065 2863 53111
rect 2941 53065 2987 53111
rect 3065 53065 3111 53111
rect 3189 53065 3235 53111
rect 3313 53065 3359 53111
rect 3437 53065 3483 53111
rect 3561 53065 3607 53111
rect 3685 53065 3731 53111
rect 3809 53065 3855 53111
rect 3933 53065 3979 53111
rect 4057 53065 4103 53111
rect 4181 53065 4227 53111
rect 4305 53065 4351 53111
rect 4429 53065 4475 53111
rect 4553 53065 4599 53111
rect 4677 53065 4723 53111
rect 4801 53065 4847 53111
rect 4925 53065 4971 53111
rect 5049 53065 5095 53111
rect 5173 53065 5219 53111
rect 5297 53065 5343 53111
rect 5421 53065 5467 53111
rect 5545 53065 5591 53111
rect 5669 53065 5715 53111
rect 5793 53065 5839 53111
rect 5917 53065 5963 53111
rect 6041 53065 6087 53111
rect 6165 53065 6211 53111
rect 6289 53065 6335 53111
rect 6413 53065 6459 53111
rect 6537 53065 6583 53111
rect 6661 53065 6707 53111
rect 6785 53065 6831 53111
rect 6909 53065 6955 53111
rect 7033 53065 7079 53111
rect 7157 53065 7203 53111
rect 7281 53065 7327 53111
rect 7405 53065 7451 53111
rect 7529 53065 7575 53111
rect 7653 53065 7699 53111
rect 7777 53065 7823 53111
rect 7901 53065 7947 53111
rect 8025 53065 8071 53111
rect 8149 53065 8195 53111
rect 8273 53065 8319 53111
rect 8397 53065 8443 53111
rect 8521 53065 8567 53111
rect 8645 53065 8691 53111
rect 8769 53065 8815 53111
rect 8893 53065 8939 53111
rect 9017 53065 9063 53111
rect 9141 53065 9187 53111
rect 9265 53065 9311 53111
rect 9389 53065 9435 53111
rect 9513 53065 9559 53111
rect 9637 53065 9683 53111
rect 9761 53065 9807 53111
rect 9885 53065 9931 53111
rect 10009 53065 10055 53111
rect 10133 53065 10179 53111
rect 10257 53065 10303 53111
rect 10381 53065 10427 53111
rect 10505 53065 10551 53111
rect 10629 53065 10675 53111
rect 10753 53065 10799 53111
rect 10877 53065 10923 53111
rect 11001 53065 11047 53111
rect 11125 53065 11171 53111
rect 11249 53065 11295 53111
rect 11373 53065 11419 53111
rect 11497 53065 11543 53111
rect 11621 53065 11667 53111
rect 11745 53065 11791 53111
rect 11869 53065 11915 53111
rect 11993 53065 12039 53111
rect 12117 53065 12163 53111
rect 12241 53065 12287 53111
rect 12365 53065 12411 53111
rect 12489 53065 12535 53111
rect 12613 53065 12659 53111
rect 12737 53065 12783 53111
rect 12861 53065 12907 53111
rect 12985 53065 13031 53111
rect 13109 53065 13155 53111
rect 13233 53065 13279 53111
rect 13357 53065 13403 53111
rect 13481 53065 13527 53111
rect 13605 53065 13651 53111
rect 13729 53065 13775 53111
rect 13853 53065 13899 53111
rect 13977 53065 14023 53111
rect 14101 53065 14147 53111
rect 14225 53065 14271 53111
rect 14349 53065 14395 53111
rect 14473 53065 14519 53111
rect 14597 53065 14643 53111
rect 14721 53065 14767 53111
rect 14845 53065 14891 53111
rect 14969 53065 15015 53111
rect 15093 53065 15139 53111
rect 15217 53065 15263 53111
rect 15341 53065 15387 53111
rect 15465 53065 15511 53111
rect 15589 53065 15635 53111
rect 15713 53065 15759 53111
rect 15837 53065 15883 53111
rect 15961 53065 16007 53111
rect 16085 53065 16131 53111
rect 16209 53065 16255 53111
rect 16333 53065 16379 53111
rect 16457 53065 16503 53111
rect 16581 53065 16627 53111
rect 16705 53065 16751 53111
rect 16829 53065 16875 53111
rect 16953 53065 16999 53111
rect 17077 53065 17123 53111
rect 17201 53065 17247 53111
rect 17325 53065 17371 53111
rect 17449 53065 17495 53111
rect 17573 53065 17619 53111
rect 17697 53065 17743 53111
rect 17821 53065 17867 53111
rect 17945 53065 17991 53111
rect 18069 53065 18115 53111
rect 18193 53065 18239 53111
rect 18317 53065 18363 53111
rect 18441 53065 18487 53111
rect 18565 53065 18611 53111
rect 18689 53065 18735 53111
rect 18813 53065 18859 53111
rect 18937 53065 18983 53111
rect 19061 53065 19107 53111
rect 19185 53065 19231 53111
rect 19309 53065 19355 53111
rect 19433 53065 19479 53111
rect 19557 53065 19603 53111
rect 19681 53065 19727 53111
rect 19805 53065 19851 53111
rect 19929 53065 19975 53111
rect 20053 53065 20099 53111
rect 20177 53065 20223 53111
rect 20301 53065 20347 53111
rect 20425 53065 20471 53111
rect 20549 53065 20595 53111
rect 20673 53065 20719 53111
rect 20797 53065 20843 53111
rect 20921 53065 20967 53111
rect 21045 53065 21091 53111
rect 21169 53065 21215 53111
rect 21293 53065 21339 53111
rect 21417 53065 21463 53111
rect 21541 53065 21587 53111
rect 21665 53065 21711 53111
rect 21789 53065 21835 53111
rect 21913 53065 21959 53111
rect 22037 53065 22083 53111
rect 22161 53065 22207 53111
rect 22285 53065 22331 53111
rect 22409 53065 22455 53111
rect 22533 53065 22579 53111
rect 22657 53065 22703 53111
rect 22781 53065 22827 53111
rect 22905 53065 22951 53111
rect 23029 53065 23075 53111
rect 23153 53065 23199 53111
rect 23277 53065 23323 53111
rect 23401 53065 23447 53111
rect 23525 53065 23571 53111
rect 23649 53065 23695 53111
rect 23773 53065 23819 53111
rect 23897 53065 23943 53111
rect 24021 53065 24067 53111
rect 24145 53065 24191 53111
rect 24269 53065 24315 53111
rect 24393 53065 24439 53111
rect 24517 53065 24563 53111
rect 24641 53065 24687 53111
rect 24765 53065 24811 53111
rect 24889 53065 24935 53111
rect 25013 53065 25059 53111
rect 25137 53065 25183 53111
rect 25261 53065 25307 53111
rect 25385 53065 25431 53111
rect 25509 53065 25555 53111
rect 25633 53065 25679 53111
rect 25757 53065 25803 53111
rect 25881 53065 25927 53111
rect 26005 53065 26051 53111
rect 26129 53065 26175 53111
rect 26253 53065 26299 53111
rect 26377 53065 26423 53111
rect 26501 53065 26547 53111
rect 26625 53065 26671 53111
rect 26749 53065 26795 53111
rect 26873 53065 26919 53111
rect 26997 53065 27043 53111
rect 27121 53065 27167 53111
rect 27245 53065 27291 53111
rect 27369 53065 27415 53111
rect 27493 53065 27539 53111
rect 27617 53065 27663 53111
rect 27741 53065 27787 53111
rect 27865 53065 27911 53111
rect 27989 53065 28035 53111
rect 28113 53065 28159 53111
rect 28237 53065 28283 53111
rect 28361 53065 28407 53111
rect 28485 53065 28531 53111
rect 28609 53065 28655 53111
rect 28733 53065 28779 53111
rect 28857 53065 28903 53111
rect 28981 53065 29027 53111
rect 29105 53065 29151 53111
rect 29229 53065 29275 53111
rect 29353 53065 29399 53111
rect 29477 53065 29523 53111
rect 29601 53065 29647 53111
rect 29725 53065 29771 53111
rect 29849 53065 29895 53111
rect 29973 53065 30019 53111
rect 30097 53065 30143 53111
rect 30221 53065 30267 53111
rect 30345 53065 30391 53111
rect 30469 53065 30515 53111
rect 30593 53065 30639 53111
rect 30717 53065 30763 53111
rect 30841 53065 30887 53111
rect 30965 53065 31011 53111
rect 31089 53065 31135 53111
rect 31213 53065 31259 53111
rect 31337 53065 31383 53111
rect 31461 53065 31507 53111
rect 31585 53065 31631 53111
rect 31709 53065 31755 53111
rect 31833 53065 31879 53111
rect 31957 53065 32003 53111
rect 32081 53065 32127 53111
rect 32205 53065 32251 53111
rect 32329 53065 32375 53111
rect 32453 53065 32499 53111
rect 32577 53065 32623 53111
rect 32701 53065 32747 53111
rect 32825 53065 32871 53111
rect 32949 53065 32995 53111
rect 33073 53065 33119 53111
rect 33197 53065 33243 53111
rect 33321 53065 33367 53111
rect 33445 53065 33491 53111
rect 33569 53065 33615 53111
rect 33693 53065 33739 53111
rect 33817 53065 33863 53111
rect 33941 53065 33987 53111
rect 34065 53065 34111 53111
rect 34189 53065 34235 53111
rect 34313 53065 34359 53111
rect 34437 53065 34483 53111
rect 34561 53065 34607 53111
rect 34685 53065 34731 53111
rect 34809 53065 34855 53111
rect 34933 53065 34979 53111
rect 35057 53065 35103 53111
rect 35181 53065 35227 53111
rect 35305 53065 35351 53111
rect 35429 53065 35475 53111
rect 35553 53065 35599 53111
rect 35677 53065 35723 53111
rect 35801 53065 35847 53111
rect 35925 53065 35971 53111
rect 36049 53065 36095 53111
rect 36173 53065 36219 53111
rect 36297 53065 36343 53111
rect 36421 53065 36467 53111
rect 36545 53065 36591 53111
rect 36669 53065 36715 53111
rect 36793 53065 36839 53111
rect 36917 53065 36963 53111
rect 37041 53065 37087 53111
rect 37165 53065 37211 53111
rect 37289 53065 37335 53111
rect 37413 53065 37459 53111
rect 37537 53065 37583 53111
rect 37661 53065 37707 53111
rect 37785 53065 37831 53111
rect 37909 53065 37955 53111
rect 38033 53065 38079 53111
rect 38157 53065 38203 53111
rect 38281 53065 38327 53111
rect 38405 53065 38451 53111
rect 38529 53065 38575 53111
rect 38653 53065 38699 53111
rect 38777 53065 38823 53111
rect 38901 53065 38947 53111
rect 39025 53065 39071 53111
rect 39149 53065 39195 53111
rect 39273 53065 39319 53111
rect 39397 53065 39443 53111
rect 39521 53065 39567 53111
rect 39645 53065 39691 53111
rect 39769 53065 39815 53111
rect 39893 53065 39939 53111
rect 40017 53065 40063 53111
rect 40141 53065 40187 53111
rect 40265 53065 40311 53111
rect 40389 53065 40435 53111
rect 40513 53065 40559 53111
rect 40637 53065 40683 53111
rect 40761 53065 40807 53111
rect 40885 53065 40931 53111
rect 41009 53065 41055 53111
rect 41133 53065 41179 53111
rect 41257 53065 41303 53111
rect 41381 53065 41427 53111
rect 41505 53065 41551 53111
rect 41629 53065 41675 53111
rect 41753 53065 41799 53111
rect 41877 53065 41923 53111
rect 42001 53065 42047 53111
rect 42125 53065 42171 53111
rect 42249 53065 42295 53111
rect 42373 53065 42419 53111
rect 42497 53065 42543 53111
rect 42621 53065 42667 53111
rect 42745 53065 42791 53111
rect 42869 53065 42915 53111
rect 42993 53065 43039 53111
rect 43117 53065 43163 53111
rect 43241 53065 43287 53111
rect 43365 53065 43411 53111
rect 43489 53065 43535 53111
rect 43613 53065 43659 53111
rect 43737 53065 43783 53111
rect 43861 53065 43907 53111
rect 43985 53065 44031 53111
rect 44109 53065 44155 53111
rect 44233 53065 44279 53111
rect 44357 53065 44403 53111
rect 44481 53065 44527 53111
rect 44605 53065 44651 53111
rect 44729 53065 44775 53111
rect 44853 53065 44899 53111
rect 44977 53065 45023 53111
rect 45101 53065 45147 53111
rect 45225 53065 45271 53111
rect 45349 53065 45395 53111
rect 45473 53065 45519 53111
rect 45597 53065 45643 53111
rect 45721 53065 45767 53111
rect 45845 53065 45891 53111
rect 45969 53065 46015 53111
rect 46093 53065 46139 53111
rect 46217 53065 46263 53111
rect 46341 53065 46387 53111
rect 46465 53065 46511 53111
rect 46589 53065 46635 53111
rect 46713 53065 46759 53111
rect 46837 53065 46883 53111
rect 46961 53065 47007 53111
rect 47085 53065 47131 53111
rect 47209 53065 47255 53111
rect 47333 53065 47379 53111
rect 47457 53065 47503 53111
rect 47581 53065 47627 53111
rect 47705 53065 47751 53111
rect 47829 53065 47875 53111
rect 47953 53065 47999 53111
rect 48077 53065 48123 53111
rect 48201 53065 48247 53111
rect 48325 53065 48371 53111
rect 48449 53065 48495 53111
rect 48573 53065 48619 53111
rect 48697 53065 48743 53111
rect 48821 53065 48867 53111
rect 48945 53065 48991 53111
rect 49069 53065 49115 53111
rect 49193 53065 49239 53111
rect 49317 53065 49363 53111
rect 49441 53065 49487 53111
rect 49565 53065 49611 53111
rect 49689 53065 49735 53111
rect 49813 53065 49859 53111
rect 49937 53065 49983 53111
rect 50061 53065 50107 53111
rect 50185 53065 50231 53111
rect 50309 53065 50355 53111
rect 50433 53065 50479 53111
rect 50557 53065 50603 53111
rect 50681 53065 50727 53111
rect 50805 53065 50851 53111
rect 50929 53065 50975 53111
rect 51053 53065 51099 53111
rect 51177 53065 51223 53111
rect 51301 53065 51347 53111
rect 51425 53065 51471 53111
rect 51549 53065 51595 53111
rect 51673 53065 51719 53111
rect 51797 53065 51843 53111
rect 51921 53065 51967 53111
rect 52045 53065 52091 53111
rect 52169 53065 52215 53111
rect 52293 53065 52339 53111
rect 52417 53065 52463 53111
rect 52541 53065 52587 53111
rect 52665 53065 52711 53111
rect 52789 53065 52835 53111
rect 52913 53065 52959 53111
rect 53037 53065 53083 53111
rect 53161 53065 53207 53111
rect 53285 53065 53331 53111
rect 53409 53065 53455 53111
rect 53533 53065 53579 53111
rect 53657 53065 53703 53111
rect 53781 53065 53827 53111
rect 53905 53065 53951 53111
rect 54029 53065 54075 53111
rect 54153 53065 54199 53111
rect 54277 53065 54323 53111
rect 54401 53065 54447 53111
rect 54525 53065 54571 53111
rect 54649 53065 54695 53111
rect 54773 53065 54819 53111
rect 54897 53065 54943 53111
rect 55021 53065 55067 53111
rect 55145 53065 55191 53111
rect 55269 53065 55315 53111
rect 55393 53065 55439 53111
rect 55517 53065 55563 53111
rect 55641 53065 55687 53111
rect 55765 53065 55811 53111
rect 55889 53065 55935 53111
rect 56013 53065 56059 53111
rect 56137 53065 56183 53111
rect 56261 53065 56307 53111
rect 56385 53065 56431 53111
rect 56509 53065 56555 53111
rect 56633 53065 56679 53111
rect 56757 53065 56803 53111
rect 56881 53065 56927 53111
rect 57005 53065 57051 53111
rect 57129 53065 57175 53111
rect 57253 53065 57299 53111
rect 57377 53065 57423 53111
rect 57501 53065 57547 53111
rect 57625 53065 57671 53111
rect 57749 53065 57795 53111
rect 57873 53065 57919 53111
rect 57997 53065 58043 53111
rect 58121 53065 58167 53111
rect 58245 53065 58291 53111
rect 58369 53065 58415 53111
rect 58493 53065 58539 53111
rect 58617 53065 58663 53111
rect 58741 53065 58787 53111
rect 58865 53065 58911 53111
rect 58989 53065 59035 53111
rect 59113 53065 59159 53111
rect 59237 53065 59283 53111
rect 59361 53065 59407 53111
rect 59485 53065 59531 53111
rect 59609 53065 59655 53111
rect 59733 53065 59779 53111
rect 59857 53065 59903 53111
rect 59981 53065 60027 53111
rect 60105 53065 60151 53111
rect 60229 53065 60275 53111
rect 60353 53065 60399 53111
rect 60477 53065 60523 53111
rect 60601 53065 60647 53111
rect 60725 53065 60771 53111
rect 60849 53065 60895 53111
rect 60973 53065 61019 53111
rect 61097 53065 61143 53111
rect 61221 53065 61267 53111
rect 61345 53065 61391 53111
rect 61469 53065 61515 53111
rect 61593 53065 61639 53111
rect 61717 53065 61763 53111
rect 61841 53065 61887 53111
rect 61965 53065 62011 53111
rect 62089 53065 62135 53111
rect 62213 53065 62259 53111
rect 62337 53065 62383 53111
rect 62461 53065 62507 53111
rect 62585 53065 62631 53111
rect 62709 53065 62755 53111
rect 62833 53065 62879 53111
rect 62957 53065 63003 53111
rect 63081 53065 63127 53111
rect 63205 53065 63251 53111
rect 63329 53065 63375 53111
rect 63453 53065 63499 53111
rect 63577 53065 63623 53111
rect 63701 53065 63747 53111
rect 63825 53065 63871 53111
rect 63949 53065 63995 53111
rect 64073 53065 64119 53111
rect 64197 53065 64243 53111
rect 64321 53065 64367 53111
rect 64445 53065 64491 53111
rect 64569 53065 64615 53111
rect 64693 53065 64739 53111
rect 64817 53065 64863 53111
rect 64941 53065 64987 53111
rect 65065 53065 65111 53111
rect 65189 53065 65235 53111
rect 65313 53065 65359 53111
rect 65437 53065 65483 53111
rect 65561 53065 65607 53111
rect 65685 53065 65731 53111
rect 65809 53065 65855 53111
rect 65933 53065 65979 53111
rect 66057 53065 66103 53111
rect 66181 53065 66227 53111
rect 66305 53065 66351 53111
rect 66429 53065 66475 53111
rect 66553 53065 66599 53111
rect 66677 53065 66723 53111
rect 66801 53065 66847 53111
rect 66925 53065 66971 53111
rect 67049 53065 67095 53111
rect 67173 53065 67219 53111
rect 67297 53065 67343 53111
rect 67421 53065 67467 53111
rect 67545 53065 67591 53111
rect 67669 53065 67715 53111
rect 67793 53065 67839 53111
rect 67917 53065 67963 53111
rect 68041 53065 68087 53111
rect 68165 53065 68211 53111
rect 68289 53065 68335 53111
rect 68413 53065 68459 53111
rect 68537 53065 68583 53111
rect 68661 53065 68707 53111
rect 68785 53065 68831 53111
rect 68909 53065 68955 53111
rect 69033 53065 69079 53111
rect 69157 53065 69203 53111
rect 69281 53065 69327 53111
rect 69405 53065 69451 53111
rect 69529 53065 69575 53111
rect 69653 53065 69699 53111
rect 69777 53065 69823 53111
rect 69901 53065 69947 53111
rect 70025 53065 70071 53111
rect 70149 53065 70195 53111
rect 70273 53065 70319 53111
rect 70397 53065 70443 53111
rect 70521 53065 70567 53111
rect 70645 53065 70691 53111
rect 70769 53065 70815 53111
rect 70893 53065 70939 53111
rect 71017 53065 71063 53111
rect 71141 53065 71187 53111
rect 71265 53065 71311 53111
rect 71389 53065 71435 53111
rect 71513 53065 71559 53111
rect 71637 53065 71683 53111
rect 71761 53065 71807 53111
rect 71885 53065 71931 53111
rect 72009 53065 72055 53111
rect 72133 53065 72179 53111
rect 72257 53065 72303 53111
rect 72381 53065 72427 53111
rect 72505 53065 72551 53111
rect 72629 53065 72675 53111
rect 72753 53065 72799 53111
rect 72877 53065 72923 53111
rect 73001 53065 73047 53111
rect 73125 53065 73171 53111
rect 73249 53065 73295 53111
rect 73373 53065 73419 53111
rect 73497 53065 73543 53111
rect 73621 53065 73667 53111
rect 73745 53065 73791 53111
rect 73869 53065 73915 53111
rect 73993 53065 74039 53111
rect 74117 53065 74163 53111
rect 74241 53065 74287 53111
rect 74365 53065 74411 53111
rect 74489 53065 74535 53111
rect 74613 53065 74659 53111
rect 74737 53065 74783 53111
rect 74861 53065 74907 53111
rect 74985 53065 75031 53111
rect 75109 53065 75155 53111
rect 75233 53065 75279 53111
rect 75357 53065 75403 53111
rect 75481 53065 75527 53111
rect 75605 53065 75651 53111
rect 75729 53065 75775 53111
rect 75853 53065 75899 53111
rect 75977 53065 76023 53111
rect 76101 53065 76147 53111
rect 76225 53065 76271 53111
rect 76349 53065 76395 53111
rect 76473 53065 76519 53111
rect 76597 53065 76643 53111
rect 76721 53065 76767 53111
rect 76845 53065 76891 53111
rect 76969 53065 77015 53111
rect 77093 53065 77139 53111
rect 77217 53065 77263 53111
rect 77341 53065 77387 53111
rect 77465 53065 77511 53111
rect 77589 53065 77635 53111
rect 77713 53065 77759 53111
rect 77837 53065 77883 53111
rect 77961 53065 78007 53111
rect 78085 53065 78131 53111
rect 78209 53065 78255 53111
rect 78333 53065 78379 53111
rect 78457 53065 78503 53111
rect 78581 53065 78627 53111
rect 78705 53065 78751 53111
rect 78829 53065 78875 53111
rect 78953 53065 78999 53111
rect 79077 53065 79123 53111
rect 79201 53065 79247 53111
rect 79325 53065 79371 53111
rect 79449 53065 79495 53111
rect 79573 53065 79619 53111
rect 79697 53065 79743 53111
rect 79821 53065 79867 53111
rect 79945 53065 79991 53111
rect 80069 53065 80115 53111
rect 80193 53065 80239 53111
rect 80317 53065 80363 53111
rect 80441 53065 80487 53111
rect 80565 53065 80611 53111
rect 80689 53065 80735 53111
rect 80813 53065 80859 53111
rect 80937 53065 80983 53111
rect 81061 53065 81107 53111
rect 81185 53065 81231 53111
rect 81309 53065 81355 53111
rect 81433 53065 81479 53111
rect 81557 53065 81603 53111
rect 81681 53065 81727 53111
rect 81805 53065 81851 53111
rect 81929 53065 81975 53111
rect 82053 53065 82099 53111
rect 82177 53065 82223 53111
rect 82301 53065 82347 53111
rect 82425 53065 82471 53111
rect 82549 53065 82595 53111
rect 82673 53065 82719 53111
rect 82797 53065 82843 53111
rect 82921 53065 82967 53111
rect 83045 53065 83091 53111
rect 83169 53065 83215 53111
rect 83293 53065 83339 53111
rect 83417 53065 83463 53111
rect 83541 53065 83587 53111
rect 83665 53065 83711 53111
rect 83789 53065 83835 53111
rect 83913 53065 83959 53111
rect 84037 53065 84083 53111
rect 84161 53065 84207 53111
rect 84285 53065 84331 53111
rect 84409 53065 84455 53111
rect 84533 53065 84579 53111
rect 84657 53065 84703 53111
rect 84781 53065 84827 53111
rect 84905 53065 84951 53111
rect 85029 53065 85075 53111
rect 85153 53065 85199 53111
rect 85277 53065 85323 53111
rect 85401 53065 85447 53111
rect 85525 53065 85571 53111
rect 85649 53065 85695 53111
rect 89 1117 435 52963
rect 85451 1117 85797 52963
rect 89 969 135 1015
rect 213 969 259 1015
rect 337 969 383 1015
rect 461 969 507 1015
rect 585 969 631 1015
rect 709 969 755 1015
rect 833 969 879 1015
rect 957 969 1003 1015
rect 1081 969 1127 1015
rect 1205 969 1251 1015
rect 1329 969 1375 1015
rect 1453 969 1499 1015
rect 1577 969 1623 1015
rect 1701 969 1747 1015
rect 1825 969 1871 1015
rect 1949 969 1995 1015
rect 2073 969 2119 1015
rect 2197 969 2243 1015
rect 2321 969 2367 1015
rect 2445 969 2491 1015
rect 2569 969 2615 1015
rect 2693 969 2739 1015
rect 2817 969 2863 1015
rect 2941 969 2987 1015
rect 3065 969 3111 1015
rect 3189 969 3235 1015
rect 3313 969 3359 1015
rect 3437 969 3483 1015
rect 3561 969 3607 1015
rect 3685 969 3731 1015
rect 3809 969 3855 1015
rect 3933 969 3979 1015
rect 4057 969 4103 1015
rect 4181 969 4227 1015
rect 4305 969 4351 1015
rect 4429 969 4475 1015
rect 4553 969 4599 1015
rect 4677 969 4723 1015
rect 4801 969 4847 1015
rect 4925 969 4971 1015
rect 5049 969 5095 1015
rect 5173 969 5219 1015
rect 5297 969 5343 1015
rect 5421 969 5467 1015
rect 5545 969 5591 1015
rect 5669 969 5715 1015
rect 5793 969 5839 1015
rect 5917 969 5963 1015
rect 6041 969 6087 1015
rect 6165 969 6211 1015
rect 6289 969 6335 1015
rect 6413 969 6459 1015
rect 6537 969 6583 1015
rect 6661 969 6707 1015
rect 6785 969 6831 1015
rect 6909 969 6955 1015
rect 7033 969 7079 1015
rect 7157 969 7203 1015
rect 7281 969 7327 1015
rect 7405 969 7451 1015
rect 7529 969 7575 1015
rect 7653 969 7699 1015
rect 7777 969 7823 1015
rect 7901 969 7947 1015
rect 8025 969 8071 1015
rect 8149 969 8195 1015
rect 8273 969 8319 1015
rect 8397 969 8443 1015
rect 8521 969 8567 1015
rect 8645 969 8691 1015
rect 8769 969 8815 1015
rect 8893 969 8939 1015
rect 9017 969 9063 1015
rect 9141 969 9187 1015
rect 9265 969 9311 1015
rect 9389 969 9435 1015
rect 9513 969 9559 1015
rect 9637 969 9683 1015
rect 9761 969 9807 1015
rect 9885 969 9931 1015
rect 10009 969 10055 1015
rect 10133 969 10179 1015
rect 10257 969 10303 1015
rect 10381 969 10427 1015
rect 10505 969 10551 1015
rect 10629 969 10675 1015
rect 10753 969 10799 1015
rect 10877 969 10923 1015
rect 11001 969 11047 1015
rect 11125 969 11171 1015
rect 11249 969 11295 1015
rect 11373 969 11419 1015
rect 11497 969 11543 1015
rect 11621 969 11667 1015
rect 11745 969 11791 1015
rect 11869 969 11915 1015
rect 11993 969 12039 1015
rect 12117 969 12163 1015
rect 12241 969 12287 1015
rect 12365 969 12411 1015
rect 12489 969 12535 1015
rect 12613 969 12659 1015
rect 12737 969 12783 1015
rect 12861 969 12907 1015
rect 12985 969 13031 1015
rect 13109 969 13155 1015
rect 13233 969 13279 1015
rect 13357 969 13403 1015
rect 13481 969 13527 1015
rect 13605 969 13651 1015
rect 13729 969 13775 1015
rect 13853 969 13899 1015
rect 13977 969 14023 1015
rect 14101 969 14147 1015
rect 14225 969 14271 1015
rect 14349 969 14395 1015
rect 14473 969 14519 1015
rect 14597 969 14643 1015
rect 14721 969 14767 1015
rect 14845 969 14891 1015
rect 14969 969 15015 1015
rect 15093 969 15139 1015
rect 15217 969 15263 1015
rect 15341 969 15387 1015
rect 15465 969 15511 1015
rect 15589 969 15635 1015
rect 15713 969 15759 1015
rect 15837 969 15883 1015
rect 15961 969 16007 1015
rect 16085 969 16131 1015
rect 16209 969 16255 1015
rect 16333 969 16379 1015
rect 16457 969 16503 1015
rect 16581 969 16627 1015
rect 16705 969 16751 1015
rect 16829 969 16875 1015
rect 16953 969 16999 1015
rect 17077 969 17123 1015
rect 17201 969 17247 1015
rect 17325 969 17371 1015
rect 17449 969 17495 1015
rect 17573 969 17619 1015
rect 17697 969 17743 1015
rect 17821 969 17867 1015
rect 17945 969 17991 1015
rect 18069 969 18115 1015
rect 18193 969 18239 1015
rect 18317 969 18363 1015
rect 18441 969 18487 1015
rect 18565 969 18611 1015
rect 18689 969 18735 1015
rect 18813 969 18859 1015
rect 18937 969 18983 1015
rect 19061 969 19107 1015
rect 19185 969 19231 1015
rect 19309 969 19355 1015
rect 19433 969 19479 1015
rect 19557 969 19603 1015
rect 19681 969 19727 1015
rect 19805 969 19851 1015
rect 19929 969 19975 1015
rect 20053 969 20099 1015
rect 20177 969 20223 1015
rect 20301 969 20347 1015
rect 20425 969 20471 1015
rect 20549 969 20595 1015
rect 20673 969 20719 1015
rect 20797 969 20843 1015
rect 20921 969 20967 1015
rect 21045 969 21091 1015
rect 21169 969 21215 1015
rect 21293 969 21339 1015
rect 21417 969 21463 1015
rect 21541 969 21587 1015
rect 21665 969 21711 1015
rect 21789 969 21835 1015
rect 21913 969 21959 1015
rect 22037 969 22083 1015
rect 22161 969 22207 1015
rect 22285 969 22331 1015
rect 22409 969 22455 1015
rect 22533 969 22579 1015
rect 22657 969 22703 1015
rect 22781 969 22827 1015
rect 22905 969 22951 1015
rect 23029 969 23075 1015
rect 23153 969 23199 1015
rect 23277 969 23323 1015
rect 23401 969 23447 1015
rect 23525 969 23571 1015
rect 23649 969 23695 1015
rect 23773 969 23819 1015
rect 23897 969 23943 1015
rect 24021 969 24067 1015
rect 24145 969 24191 1015
rect 24269 969 24315 1015
rect 24393 969 24439 1015
rect 24517 969 24563 1015
rect 24641 969 24687 1015
rect 24765 969 24811 1015
rect 24889 969 24935 1015
rect 25013 969 25059 1015
rect 25137 969 25183 1015
rect 25261 969 25307 1015
rect 25385 969 25431 1015
rect 25509 969 25555 1015
rect 25633 969 25679 1015
rect 25757 969 25803 1015
rect 25881 969 25927 1015
rect 26005 969 26051 1015
rect 26129 969 26175 1015
rect 26253 969 26299 1015
rect 26377 969 26423 1015
rect 26501 969 26547 1015
rect 26625 969 26671 1015
rect 26749 969 26795 1015
rect 26873 969 26919 1015
rect 26997 969 27043 1015
rect 27121 969 27167 1015
rect 27245 969 27291 1015
rect 27369 969 27415 1015
rect 27493 969 27539 1015
rect 27617 969 27663 1015
rect 27741 969 27787 1015
rect 27865 969 27911 1015
rect 27989 969 28035 1015
rect 28113 969 28159 1015
rect 28237 969 28283 1015
rect 28361 969 28407 1015
rect 28485 969 28531 1015
rect 28609 969 28655 1015
rect 28733 969 28779 1015
rect 28857 969 28903 1015
rect 28981 969 29027 1015
rect 29105 969 29151 1015
rect 29229 969 29275 1015
rect 29353 969 29399 1015
rect 29477 969 29523 1015
rect 29601 969 29647 1015
rect 29725 969 29771 1015
rect 29849 969 29895 1015
rect 29973 969 30019 1015
rect 30097 969 30143 1015
rect 30221 969 30267 1015
rect 30345 969 30391 1015
rect 30469 969 30515 1015
rect 30593 969 30639 1015
rect 30717 969 30763 1015
rect 30841 969 30887 1015
rect 30965 969 31011 1015
rect 31089 969 31135 1015
rect 31213 969 31259 1015
rect 31337 969 31383 1015
rect 31461 969 31507 1015
rect 31585 969 31631 1015
rect 31709 969 31755 1015
rect 31833 969 31879 1015
rect 31957 969 32003 1015
rect 32081 969 32127 1015
rect 32205 969 32251 1015
rect 32329 969 32375 1015
rect 32453 969 32499 1015
rect 32577 969 32623 1015
rect 32701 969 32747 1015
rect 32825 969 32871 1015
rect 32949 969 32995 1015
rect 33073 969 33119 1015
rect 33197 969 33243 1015
rect 33321 969 33367 1015
rect 33445 969 33491 1015
rect 33569 969 33615 1015
rect 33693 969 33739 1015
rect 33817 969 33863 1015
rect 33941 969 33987 1015
rect 34065 969 34111 1015
rect 34189 969 34235 1015
rect 34313 969 34359 1015
rect 34437 969 34483 1015
rect 34561 969 34607 1015
rect 34685 969 34731 1015
rect 34809 969 34855 1015
rect 34933 969 34979 1015
rect 35057 969 35103 1015
rect 35181 969 35227 1015
rect 35305 969 35351 1015
rect 35429 969 35475 1015
rect 35553 969 35599 1015
rect 35677 969 35723 1015
rect 35801 969 35847 1015
rect 35925 969 35971 1015
rect 36049 969 36095 1015
rect 36173 969 36219 1015
rect 36297 969 36343 1015
rect 36421 969 36467 1015
rect 36545 969 36591 1015
rect 36669 969 36715 1015
rect 36793 969 36839 1015
rect 36917 969 36963 1015
rect 37041 969 37087 1015
rect 37165 969 37211 1015
rect 37289 969 37335 1015
rect 37413 969 37459 1015
rect 37537 969 37583 1015
rect 37661 969 37707 1015
rect 37785 969 37831 1015
rect 37909 969 37955 1015
rect 38033 969 38079 1015
rect 38157 969 38203 1015
rect 38281 969 38327 1015
rect 38405 969 38451 1015
rect 38529 969 38575 1015
rect 38653 969 38699 1015
rect 38777 969 38823 1015
rect 38901 969 38947 1015
rect 39025 969 39071 1015
rect 39149 969 39195 1015
rect 39273 969 39319 1015
rect 39397 969 39443 1015
rect 39521 969 39567 1015
rect 39645 969 39691 1015
rect 39769 969 39815 1015
rect 39893 969 39939 1015
rect 40017 969 40063 1015
rect 40141 969 40187 1015
rect 40265 969 40311 1015
rect 40389 969 40435 1015
rect 40513 969 40559 1015
rect 40637 969 40683 1015
rect 40761 969 40807 1015
rect 40885 969 40931 1015
rect 41009 969 41055 1015
rect 41133 969 41179 1015
rect 41257 969 41303 1015
rect 41381 969 41427 1015
rect 41505 969 41551 1015
rect 41629 969 41675 1015
rect 41753 969 41799 1015
rect 41877 969 41923 1015
rect 42001 969 42047 1015
rect 42125 969 42171 1015
rect 42249 969 42295 1015
rect 42373 969 42419 1015
rect 42497 969 42543 1015
rect 42621 969 42667 1015
rect 42745 969 42791 1015
rect 42869 969 42915 1015
rect 42993 969 43039 1015
rect 43117 969 43163 1015
rect 43241 969 43287 1015
rect 43365 969 43411 1015
rect 43489 969 43535 1015
rect 43613 969 43659 1015
rect 43737 969 43783 1015
rect 43861 969 43907 1015
rect 43985 969 44031 1015
rect 44109 969 44155 1015
rect 44233 969 44279 1015
rect 44357 969 44403 1015
rect 44481 969 44527 1015
rect 44605 969 44651 1015
rect 44729 969 44775 1015
rect 44853 969 44899 1015
rect 44977 969 45023 1015
rect 45101 969 45147 1015
rect 45225 969 45271 1015
rect 45349 969 45395 1015
rect 45473 969 45519 1015
rect 45597 969 45643 1015
rect 45721 969 45767 1015
rect 45845 969 45891 1015
rect 45969 969 46015 1015
rect 46093 969 46139 1015
rect 46217 969 46263 1015
rect 46341 969 46387 1015
rect 46465 969 46511 1015
rect 46589 969 46635 1015
rect 46713 969 46759 1015
rect 46837 969 46883 1015
rect 46961 969 47007 1015
rect 47085 969 47131 1015
rect 47209 969 47255 1015
rect 47333 969 47379 1015
rect 47457 969 47503 1015
rect 47581 969 47627 1015
rect 47705 969 47751 1015
rect 47829 969 47875 1015
rect 47953 969 47999 1015
rect 48077 969 48123 1015
rect 48201 969 48247 1015
rect 48325 969 48371 1015
rect 48449 969 48495 1015
rect 48573 969 48619 1015
rect 48697 969 48743 1015
rect 48821 969 48867 1015
rect 48945 969 48991 1015
rect 49069 969 49115 1015
rect 49193 969 49239 1015
rect 49317 969 49363 1015
rect 49441 969 49487 1015
rect 49565 969 49611 1015
rect 49689 969 49735 1015
rect 49813 969 49859 1015
rect 49937 969 49983 1015
rect 50061 969 50107 1015
rect 50185 969 50231 1015
rect 50309 969 50355 1015
rect 50433 969 50479 1015
rect 50557 969 50603 1015
rect 50681 969 50727 1015
rect 50805 969 50851 1015
rect 50929 969 50975 1015
rect 51053 969 51099 1015
rect 51177 969 51223 1015
rect 51301 969 51347 1015
rect 51425 969 51471 1015
rect 51549 969 51595 1015
rect 51673 969 51719 1015
rect 51797 969 51843 1015
rect 51921 969 51967 1015
rect 52045 969 52091 1015
rect 52169 969 52215 1015
rect 52293 969 52339 1015
rect 52417 969 52463 1015
rect 52541 969 52587 1015
rect 52665 969 52711 1015
rect 52789 969 52835 1015
rect 52913 969 52959 1015
rect 53037 969 53083 1015
rect 53161 969 53207 1015
rect 53285 969 53331 1015
rect 53409 969 53455 1015
rect 53533 969 53579 1015
rect 53657 969 53703 1015
rect 53781 969 53827 1015
rect 53905 969 53951 1015
rect 54029 969 54075 1015
rect 54153 969 54199 1015
rect 54277 969 54323 1015
rect 54401 969 54447 1015
rect 54525 969 54571 1015
rect 54649 969 54695 1015
rect 54773 969 54819 1015
rect 54897 969 54943 1015
rect 55021 969 55067 1015
rect 55145 969 55191 1015
rect 55269 969 55315 1015
rect 55393 969 55439 1015
rect 55517 969 55563 1015
rect 55641 969 55687 1015
rect 55765 969 55811 1015
rect 55889 969 55935 1015
rect 56013 969 56059 1015
rect 56137 969 56183 1015
rect 56261 969 56307 1015
rect 56385 969 56431 1015
rect 56509 969 56555 1015
rect 56633 969 56679 1015
rect 56757 969 56803 1015
rect 56881 969 56927 1015
rect 57005 969 57051 1015
rect 57129 969 57175 1015
rect 57253 969 57299 1015
rect 57377 969 57423 1015
rect 57501 969 57547 1015
rect 57625 969 57671 1015
rect 57749 969 57795 1015
rect 57873 969 57919 1015
rect 57997 969 58043 1015
rect 58121 969 58167 1015
rect 58245 969 58291 1015
rect 58369 969 58415 1015
rect 58493 969 58539 1015
rect 58617 969 58663 1015
rect 58741 969 58787 1015
rect 58865 969 58911 1015
rect 58989 969 59035 1015
rect 59113 969 59159 1015
rect 59237 969 59283 1015
rect 59361 969 59407 1015
rect 59485 969 59531 1015
rect 59609 969 59655 1015
rect 59733 969 59779 1015
rect 59857 969 59903 1015
rect 59981 969 60027 1015
rect 60105 969 60151 1015
rect 60229 969 60275 1015
rect 60353 969 60399 1015
rect 60477 969 60523 1015
rect 60601 969 60647 1015
rect 60725 969 60771 1015
rect 60849 969 60895 1015
rect 60973 969 61019 1015
rect 61097 969 61143 1015
rect 61221 969 61267 1015
rect 61345 969 61391 1015
rect 61469 969 61515 1015
rect 61593 969 61639 1015
rect 61717 969 61763 1015
rect 61841 969 61887 1015
rect 61965 969 62011 1015
rect 62089 969 62135 1015
rect 62213 969 62259 1015
rect 62337 969 62383 1015
rect 62461 969 62507 1015
rect 62585 969 62631 1015
rect 62709 969 62755 1015
rect 62833 969 62879 1015
rect 62957 969 63003 1015
rect 63081 969 63127 1015
rect 63205 969 63251 1015
rect 63329 969 63375 1015
rect 63453 969 63499 1015
rect 63577 969 63623 1015
rect 63701 969 63747 1015
rect 63825 969 63871 1015
rect 63949 969 63995 1015
rect 64073 969 64119 1015
rect 64197 969 64243 1015
rect 64321 969 64367 1015
rect 64445 969 64491 1015
rect 64569 969 64615 1015
rect 64693 969 64739 1015
rect 64817 969 64863 1015
rect 64941 969 64987 1015
rect 65065 969 65111 1015
rect 65189 969 65235 1015
rect 65313 969 65359 1015
rect 65437 969 65483 1015
rect 65561 969 65607 1015
rect 65685 969 65731 1015
rect 65809 969 65855 1015
rect 65933 969 65979 1015
rect 66057 969 66103 1015
rect 66181 969 66227 1015
rect 66305 969 66351 1015
rect 66429 969 66475 1015
rect 66553 969 66599 1015
rect 66677 969 66723 1015
rect 66801 969 66847 1015
rect 66925 969 66971 1015
rect 67049 969 67095 1015
rect 67173 969 67219 1015
rect 67297 969 67343 1015
rect 67421 969 67467 1015
rect 67545 969 67591 1015
rect 67669 969 67715 1015
rect 67793 969 67839 1015
rect 67917 969 67963 1015
rect 68041 969 68087 1015
rect 68165 969 68211 1015
rect 68289 969 68335 1015
rect 68413 969 68459 1015
rect 68537 969 68583 1015
rect 68661 969 68707 1015
rect 68785 969 68831 1015
rect 68909 969 68955 1015
rect 69033 969 69079 1015
rect 69157 969 69203 1015
rect 69281 969 69327 1015
rect 69405 969 69451 1015
rect 69529 969 69575 1015
rect 69653 969 69699 1015
rect 69777 969 69823 1015
rect 69901 969 69947 1015
rect 70025 969 70071 1015
rect 70149 969 70195 1015
rect 70273 969 70319 1015
rect 70397 969 70443 1015
rect 70521 969 70567 1015
rect 70645 969 70691 1015
rect 70769 969 70815 1015
rect 70893 969 70939 1015
rect 71017 969 71063 1015
rect 71141 969 71187 1015
rect 71265 969 71311 1015
rect 71389 969 71435 1015
rect 71513 969 71559 1015
rect 71637 969 71683 1015
rect 71761 969 71807 1015
rect 71885 969 71931 1015
rect 72009 969 72055 1015
rect 72133 969 72179 1015
rect 72257 969 72303 1015
rect 72381 969 72427 1015
rect 72505 969 72551 1015
rect 72629 969 72675 1015
rect 72753 969 72799 1015
rect 72877 969 72923 1015
rect 73001 969 73047 1015
rect 73125 969 73171 1015
rect 73249 969 73295 1015
rect 73373 969 73419 1015
rect 73497 969 73543 1015
rect 73621 969 73667 1015
rect 73745 969 73791 1015
rect 73869 969 73915 1015
rect 73993 969 74039 1015
rect 74117 969 74163 1015
rect 74241 969 74287 1015
rect 74365 969 74411 1015
rect 74489 969 74535 1015
rect 74613 969 74659 1015
rect 74737 969 74783 1015
rect 74861 969 74907 1015
rect 74985 969 75031 1015
rect 75109 969 75155 1015
rect 75233 969 75279 1015
rect 75357 969 75403 1015
rect 75481 969 75527 1015
rect 75605 969 75651 1015
rect 75729 969 75775 1015
rect 75853 969 75899 1015
rect 75977 969 76023 1015
rect 76101 969 76147 1015
rect 76225 969 76271 1015
rect 76349 969 76395 1015
rect 76473 969 76519 1015
rect 76597 969 76643 1015
rect 76721 969 76767 1015
rect 76845 969 76891 1015
rect 76969 969 77015 1015
rect 77093 969 77139 1015
rect 77217 969 77263 1015
rect 77341 969 77387 1015
rect 77465 969 77511 1015
rect 77589 969 77635 1015
rect 77713 969 77759 1015
rect 77837 969 77883 1015
rect 77961 969 78007 1015
rect 78085 969 78131 1015
rect 78209 969 78255 1015
rect 78333 969 78379 1015
rect 78457 969 78503 1015
rect 78581 969 78627 1015
rect 78705 969 78751 1015
rect 78829 969 78875 1015
rect 78953 969 78999 1015
rect 79077 969 79123 1015
rect 79201 969 79247 1015
rect 79325 969 79371 1015
rect 79449 969 79495 1015
rect 79573 969 79619 1015
rect 79697 969 79743 1015
rect 79821 969 79867 1015
rect 79945 969 79991 1015
rect 80069 969 80115 1015
rect 80193 969 80239 1015
rect 80317 969 80363 1015
rect 80441 969 80487 1015
rect 80565 969 80611 1015
rect 80689 969 80735 1015
rect 80813 969 80859 1015
rect 80937 969 80983 1015
rect 81061 969 81107 1015
rect 81185 969 81231 1015
rect 81309 969 81355 1015
rect 81433 969 81479 1015
rect 81557 969 81603 1015
rect 81681 969 81727 1015
rect 81805 969 81851 1015
rect 81929 969 81975 1015
rect 82053 969 82099 1015
rect 82177 969 82223 1015
rect 82301 969 82347 1015
rect 82425 969 82471 1015
rect 82549 969 82595 1015
rect 82673 969 82719 1015
rect 82797 969 82843 1015
rect 82921 969 82967 1015
rect 83045 969 83091 1015
rect 83169 969 83215 1015
rect 83293 969 83339 1015
rect 83417 969 83463 1015
rect 83541 969 83587 1015
rect 83665 969 83711 1015
rect 83789 969 83835 1015
rect 83913 969 83959 1015
rect 84037 969 84083 1015
rect 84161 969 84207 1015
rect 84285 969 84331 1015
rect 84409 969 84455 1015
rect 84533 969 84579 1015
rect 84657 969 84703 1015
rect 84781 969 84827 1015
rect 84905 969 84951 1015
rect 85029 969 85075 1015
rect 85153 969 85199 1015
rect 85277 969 85323 1015
rect 85401 969 85447 1015
rect 85525 969 85571 1015
rect 85649 969 85695 1015
rect 89 845 135 891
rect 213 845 259 891
rect 337 845 383 891
rect 461 845 507 891
rect 585 845 631 891
rect 709 845 755 891
rect 833 845 879 891
rect 957 845 1003 891
rect 1081 845 1127 891
rect 1205 845 1251 891
rect 1329 845 1375 891
rect 1453 845 1499 891
rect 1577 845 1623 891
rect 1701 845 1747 891
rect 1825 845 1871 891
rect 1949 845 1995 891
rect 2073 845 2119 891
rect 2197 845 2243 891
rect 2321 845 2367 891
rect 2445 845 2491 891
rect 2569 845 2615 891
rect 2693 845 2739 891
rect 2817 845 2863 891
rect 2941 845 2987 891
rect 3065 845 3111 891
rect 3189 845 3235 891
rect 3313 845 3359 891
rect 3437 845 3483 891
rect 3561 845 3607 891
rect 3685 845 3731 891
rect 3809 845 3855 891
rect 3933 845 3979 891
rect 4057 845 4103 891
rect 4181 845 4227 891
rect 4305 845 4351 891
rect 4429 845 4475 891
rect 4553 845 4599 891
rect 4677 845 4723 891
rect 4801 845 4847 891
rect 4925 845 4971 891
rect 5049 845 5095 891
rect 5173 845 5219 891
rect 5297 845 5343 891
rect 5421 845 5467 891
rect 5545 845 5591 891
rect 5669 845 5715 891
rect 5793 845 5839 891
rect 5917 845 5963 891
rect 6041 845 6087 891
rect 6165 845 6211 891
rect 6289 845 6335 891
rect 6413 845 6459 891
rect 6537 845 6583 891
rect 6661 845 6707 891
rect 6785 845 6831 891
rect 6909 845 6955 891
rect 7033 845 7079 891
rect 7157 845 7203 891
rect 7281 845 7327 891
rect 7405 845 7451 891
rect 7529 845 7575 891
rect 7653 845 7699 891
rect 7777 845 7823 891
rect 7901 845 7947 891
rect 8025 845 8071 891
rect 8149 845 8195 891
rect 8273 845 8319 891
rect 8397 845 8443 891
rect 8521 845 8567 891
rect 8645 845 8691 891
rect 8769 845 8815 891
rect 8893 845 8939 891
rect 9017 845 9063 891
rect 9141 845 9187 891
rect 9265 845 9311 891
rect 9389 845 9435 891
rect 9513 845 9559 891
rect 9637 845 9683 891
rect 9761 845 9807 891
rect 9885 845 9931 891
rect 10009 845 10055 891
rect 10133 845 10179 891
rect 10257 845 10303 891
rect 10381 845 10427 891
rect 10505 845 10551 891
rect 10629 845 10675 891
rect 10753 845 10799 891
rect 10877 845 10923 891
rect 11001 845 11047 891
rect 11125 845 11171 891
rect 11249 845 11295 891
rect 11373 845 11419 891
rect 11497 845 11543 891
rect 11621 845 11667 891
rect 11745 845 11791 891
rect 11869 845 11915 891
rect 11993 845 12039 891
rect 12117 845 12163 891
rect 12241 845 12287 891
rect 12365 845 12411 891
rect 12489 845 12535 891
rect 12613 845 12659 891
rect 12737 845 12783 891
rect 12861 845 12907 891
rect 12985 845 13031 891
rect 13109 845 13155 891
rect 13233 845 13279 891
rect 13357 845 13403 891
rect 13481 845 13527 891
rect 13605 845 13651 891
rect 13729 845 13775 891
rect 13853 845 13899 891
rect 13977 845 14023 891
rect 14101 845 14147 891
rect 14225 845 14271 891
rect 14349 845 14395 891
rect 14473 845 14519 891
rect 14597 845 14643 891
rect 14721 845 14767 891
rect 14845 845 14891 891
rect 14969 845 15015 891
rect 15093 845 15139 891
rect 15217 845 15263 891
rect 15341 845 15387 891
rect 15465 845 15511 891
rect 15589 845 15635 891
rect 15713 845 15759 891
rect 15837 845 15883 891
rect 15961 845 16007 891
rect 16085 845 16131 891
rect 16209 845 16255 891
rect 16333 845 16379 891
rect 16457 845 16503 891
rect 16581 845 16627 891
rect 16705 845 16751 891
rect 16829 845 16875 891
rect 16953 845 16999 891
rect 17077 845 17123 891
rect 17201 845 17247 891
rect 17325 845 17371 891
rect 17449 845 17495 891
rect 17573 845 17619 891
rect 17697 845 17743 891
rect 17821 845 17867 891
rect 17945 845 17991 891
rect 18069 845 18115 891
rect 18193 845 18239 891
rect 18317 845 18363 891
rect 18441 845 18487 891
rect 18565 845 18611 891
rect 18689 845 18735 891
rect 18813 845 18859 891
rect 18937 845 18983 891
rect 19061 845 19107 891
rect 19185 845 19231 891
rect 19309 845 19355 891
rect 19433 845 19479 891
rect 19557 845 19603 891
rect 19681 845 19727 891
rect 19805 845 19851 891
rect 19929 845 19975 891
rect 20053 845 20099 891
rect 20177 845 20223 891
rect 20301 845 20347 891
rect 20425 845 20471 891
rect 20549 845 20595 891
rect 20673 845 20719 891
rect 20797 845 20843 891
rect 20921 845 20967 891
rect 21045 845 21091 891
rect 21169 845 21215 891
rect 21293 845 21339 891
rect 21417 845 21463 891
rect 21541 845 21587 891
rect 21665 845 21711 891
rect 21789 845 21835 891
rect 21913 845 21959 891
rect 22037 845 22083 891
rect 22161 845 22207 891
rect 22285 845 22331 891
rect 22409 845 22455 891
rect 22533 845 22579 891
rect 22657 845 22703 891
rect 22781 845 22827 891
rect 22905 845 22951 891
rect 23029 845 23075 891
rect 23153 845 23199 891
rect 23277 845 23323 891
rect 23401 845 23447 891
rect 23525 845 23571 891
rect 23649 845 23695 891
rect 23773 845 23819 891
rect 23897 845 23943 891
rect 24021 845 24067 891
rect 24145 845 24191 891
rect 24269 845 24315 891
rect 24393 845 24439 891
rect 24517 845 24563 891
rect 24641 845 24687 891
rect 24765 845 24811 891
rect 24889 845 24935 891
rect 25013 845 25059 891
rect 25137 845 25183 891
rect 25261 845 25307 891
rect 25385 845 25431 891
rect 25509 845 25555 891
rect 25633 845 25679 891
rect 25757 845 25803 891
rect 25881 845 25927 891
rect 26005 845 26051 891
rect 26129 845 26175 891
rect 26253 845 26299 891
rect 26377 845 26423 891
rect 26501 845 26547 891
rect 26625 845 26671 891
rect 26749 845 26795 891
rect 26873 845 26919 891
rect 26997 845 27043 891
rect 27121 845 27167 891
rect 27245 845 27291 891
rect 27369 845 27415 891
rect 27493 845 27539 891
rect 27617 845 27663 891
rect 27741 845 27787 891
rect 27865 845 27911 891
rect 27989 845 28035 891
rect 28113 845 28159 891
rect 28237 845 28283 891
rect 28361 845 28407 891
rect 28485 845 28531 891
rect 28609 845 28655 891
rect 28733 845 28779 891
rect 28857 845 28903 891
rect 28981 845 29027 891
rect 29105 845 29151 891
rect 29229 845 29275 891
rect 29353 845 29399 891
rect 29477 845 29523 891
rect 29601 845 29647 891
rect 29725 845 29771 891
rect 29849 845 29895 891
rect 29973 845 30019 891
rect 30097 845 30143 891
rect 30221 845 30267 891
rect 30345 845 30391 891
rect 30469 845 30515 891
rect 30593 845 30639 891
rect 30717 845 30763 891
rect 30841 845 30887 891
rect 30965 845 31011 891
rect 31089 845 31135 891
rect 31213 845 31259 891
rect 31337 845 31383 891
rect 31461 845 31507 891
rect 31585 845 31631 891
rect 31709 845 31755 891
rect 31833 845 31879 891
rect 31957 845 32003 891
rect 32081 845 32127 891
rect 32205 845 32251 891
rect 32329 845 32375 891
rect 32453 845 32499 891
rect 32577 845 32623 891
rect 32701 845 32747 891
rect 32825 845 32871 891
rect 32949 845 32995 891
rect 33073 845 33119 891
rect 33197 845 33243 891
rect 33321 845 33367 891
rect 33445 845 33491 891
rect 33569 845 33615 891
rect 33693 845 33739 891
rect 33817 845 33863 891
rect 33941 845 33987 891
rect 34065 845 34111 891
rect 34189 845 34235 891
rect 34313 845 34359 891
rect 34437 845 34483 891
rect 34561 845 34607 891
rect 34685 845 34731 891
rect 34809 845 34855 891
rect 34933 845 34979 891
rect 35057 845 35103 891
rect 35181 845 35227 891
rect 35305 845 35351 891
rect 35429 845 35475 891
rect 35553 845 35599 891
rect 35677 845 35723 891
rect 35801 845 35847 891
rect 35925 845 35971 891
rect 36049 845 36095 891
rect 36173 845 36219 891
rect 36297 845 36343 891
rect 36421 845 36467 891
rect 36545 845 36591 891
rect 36669 845 36715 891
rect 36793 845 36839 891
rect 36917 845 36963 891
rect 37041 845 37087 891
rect 37165 845 37211 891
rect 37289 845 37335 891
rect 37413 845 37459 891
rect 37537 845 37583 891
rect 37661 845 37707 891
rect 37785 845 37831 891
rect 37909 845 37955 891
rect 38033 845 38079 891
rect 38157 845 38203 891
rect 38281 845 38327 891
rect 38405 845 38451 891
rect 38529 845 38575 891
rect 38653 845 38699 891
rect 38777 845 38823 891
rect 38901 845 38947 891
rect 39025 845 39071 891
rect 39149 845 39195 891
rect 39273 845 39319 891
rect 39397 845 39443 891
rect 39521 845 39567 891
rect 39645 845 39691 891
rect 39769 845 39815 891
rect 39893 845 39939 891
rect 40017 845 40063 891
rect 40141 845 40187 891
rect 40265 845 40311 891
rect 40389 845 40435 891
rect 40513 845 40559 891
rect 40637 845 40683 891
rect 40761 845 40807 891
rect 40885 845 40931 891
rect 41009 845 41055 891
rect 41133 845 41179 891
rect 41257 845 41303 891
rect 41381 845 41427 891
rect 41505 845 41551 891
rect 41629 845 41675 891
rect 41753 845 41799 891
rect 41877 845 41923 891
rect 42001 845 42047 891
rect 42125 845 42171 891
rect 42249 845 42295 891
rect 42373 845 42419 891
rect 42497 845 42543 891
rect 42621 845 42667 891
rect 42745 845 42791 891
rect 42869 845 42915 891
rect 42993 845 43039 891
rect 43117 845 43163 891
rect 43241 845 43287 891
rect 43365 845 43411 891
rect 43489 845 43535 891
rect 43613 845 43659 891
rect 43737 845 43783 891
rect 43861 845 43907 891
rect 43985 845 44031 891
rect 44109 845 44155 891
rect 44233 845 44279 891
rect 44357 845 44403 891
rect 44481 845 44527 891
rect 44605 845 44651 891
rect 44729 845 44775 891
rect 44853 845 44899 891
rect 44977 845 45023 891
rect 45101 845 45147 891
rect 45225 845 45271 891
rect 45349 845 45395 891
rect 45473 845 45519 891
rect 45597 845 45643 891
rect 45721 845 45767 891
rect 45845 845 45891 891
rect 45969 845 46015 891
rect 46093 845 46139 891
rect 46217 845 46263 891
rect 46341 845 46387 891
rect 46465 845 46511 891
rect 46589 845 46635 891
rect 46713 845 46759 891
rect 46837 845 46883 891
rect 46961 845 47007 891
rect 47085 845 47131 891
rect 47209 845 47255 891
rect 47333 845 47379 891
rect 47457 845 47503 891
rect 47581 845 47627 891
rect 47705 845 47751 891
rect 47829 845 47875 891
rect 47953 845 47999 891
rect 48077 845 48123 891
rect 48201 845 48247 891
rect 48325 845 48371 891
rect 48449 845 48495 891
rect 48573 845 48619 891
rect 48697 845 48743 891
rect 48821 845 48867 891
rect 48945 845 48991 891
rect 49069 845 49115 891
rect 49193 845 49239 891
rect 49317 845 49363 891
rect 49441 845 49487 891
rect 49565 845 49611 891
rect 49689 845 49735 891
rect 49813 845 49859 891
rect 49937 845 49983 891
rect 50061 845 50107 891
rect 50185 845 50231 891
rect 50309 845 50355 891
rect 50433 845 50479 891
rect 50557 845 50603 891
rect 50681 845 50727 891
rect 50805 845 50851 891
rect 50929 845 50975 891
rect 51053 845 51099 891
rect 51177 845 51223 891
rect 51301 845 51347 891
rect 51425 845 51471 891
rect 51549 845 51595 891
rect 51673 845 51719 891
rect 51797 845 51843 891
rect 51921 845 51967 891
rect 52045 845 52091 891
rect 52169 845 52215 891
rect 52293 845 52339 891
rect 52417 845 52463 891
rect 52541 845 52587 891
rect 52665 845 52711 891
rect 52789 845 52835 891
rect 52913 845 52959 891
rect 53037 845 53083 891
rect 53161 845 53207 891
rect 53285 845 53331 891
rect 53409 845 53455 891
rect 53533 845 53579 891
rect 53657 845 53703 891
rect 53781 845 53827 891
rect 53905 845 53951 891
rect 54029 845 54075 891
rect 54153 845 54199 891
rect 54277 845 54323 891
rect 54401 845 54447 891
rect 54525 845 54571 891
rect 54649 845 54695 891
rect 54773 845 54819 891
rect 54897 845 54943 891
rect 55021 845 55067 891
rect 55145 845 55191 891
rect 55269 845 55315 891
rect 55393 845 55439 891
rect 55517 845 55563 891
rect 55641 845 55687 891
rect 55765 845 55811 891
rect 55889 845 55935 891
rect 56013 845 56059 891
rect 56137 845 56183 891
rect 56261 845 56307 891
rect 56385 845 56431 891
rect 56509 845 56555 891
rect 56633 845 56679 891
rect 56757 845 56803 891
rect 56881 845 56927 891
rect 57005 845 57051 891
rect 57129 845 57175 891
rect 57253 845 57299 891
rect 57377 845 57423 891
rect 57501 845 57547 891
rect 57625 845 57671 891
rect 57749 845 57795 891
rect 57873 845 57919 891
rect 57997 845 58043 891
rect 58121 845 58167 891
rect 58245 845 58291 891
rect 58369 845 58415 891
rect 58493 845 58539 891
rect 58617 845 58663 891
rect 58741 845 58787 891
rect 58865 845 58911 891
rect 58989 845 59035 891
rect 59113 845 59159 891
rect 59237 845 59283 891
rect 59361 845 59407 891
rect 59485 845 59531 891
rect 59609 845 59655 891
rect 59733 845 59779 891
rect 59857 845 59903 891
rect 59981 845 60027 891
rect 60105 845 60151 891
rect 60229 845 60275 891
rect 60353 845 60399 891
rect 60477 845 60523 891
rect 60601 845 60647 891
rect 60725 845 60771 891
rect 60849 845 60895 891
rect 60973 845 61019 891
rect 61097 845 61143 891
rect 61221 845 61267 891
rect 61345 845 61391 891
rect 61469 845 61515 891
rect 61593 845 61639 891
rect 61717 845 61763 891
rect 61841 845 61887 891
rect 61965 845 62011 891
rect 62089 845 62135 891
rect 62213 845 62259 891
rect 62337 845 62383 891
rect 62461 845 62507 891
rect 62585 845 62631 891
rect 62709 845 62755 891
rect 62833 845 62879 891
rect 62957 845 63003 891
rect 63081 845 63127 891
rect 63205 845 63251 891
rect 63329 845 63375 891
rect 63453 845 63499 891
rect 63577 845 63623 891
rect 63701 845 63747 891
rect 63825 845 63871 891
rect 63949 845 63995 891
rect 64073 845 64119 891
rect 64197 845 64243 891
rect 64321 845 64367 891
rect 64445 845 64491 891
rect 64569 845 64615 891
rect 64693 845 64739 891
rect 64817 845 64863 891
rect 64941 845 64987 891
rect 65065 845 65111 891
rect 65189 845 65235 891
rect 65313 845 65359 891
rect 65437 845 65483 891
rect 65561 845 65607 891
rect 65685 845 65731 891
rect 65809 845 65855 891
rect 65933 845 65979 891
rect 66057 845 66103 891
rect 66181 845 66227 891
rect 66305 845 66351 891
rect 66429 845 66475 891
rect 66553 845 66599 891
rect 66677 845 66723 891
rect 66801 845 66847 891
rect 66925 845 66971 891
rect 67049 845 67095 891
rect 67173 845 67219 891
rect 67297 845 67343 891
rect 67421 845 67467 891
rect 67545 845 67591 891
rect 67669 845 67715 891
rect 67793 845 67839 891
rect 67917 845 67963 891
rect 68041 845 68087 891
rect 68165 845 68211 891
rect 68289 845 68335 891
rect 68413 845 68459 891
rect 68537 845 68583 891
rect 68661 845 68707 891
rect 68785 845 68831 891
rect 68909 845 68955 891
rect 69033 845 69079 891
rect 69157 845 69203 891
rect 69281 845 69327 891
rect 69405 845 69451 891
rect 69529 845 69575 891
rect 69653 845 69699 891
rect 69777 845 69823 891
rect 69901 845 69947 891
rect 70025 845 70071 891
rect 70149 845 70195 891
rect 70273 845 70319 891
rect 70397 845 70443 891
rect 70521 845 70567 891
rect 70645 845 70691 891
rect 70769 845 70815 891
rect 70893 845 70939 891
rect 71017 845 71063 891
rect 71141 845 71187 891
rect 71265 845 71311 891
rect 71389 845 71435 891
rect 71513 845 71559 891
rect 71637 845 71683 891
rect 71761 845 71807 891
rect 71885 845 71931 891
rect 72009 845 72055 891
rect 72133 845 72179 891
rect 72257 845 72303 891
rect 72381 845 72427 891
rect 72505 845 72551 891
rect 72629 845 72675 891
rect 72753 845 72799 891
rect 72877 845 72923 891
rect 73001 845 73047 891
rect 73125 845 73171 891
rect 73249 845 73295 891
rect 73373 845 73419 891
rect 73497 845 73543 891
rect 73621 845 73667 891
rect 73745 845 73791 891
rect 73869 845 73915 891
rect 73993 845 74039 891
rect 74117 845 74163 891
rect 74241 845 74287 891
rect 74365 845 74411 891
rect 74489 845 74535 891
rect 74613 845 74659 891
rect 74737 845 74783 891
rect 74861 845 74907 891
rect 74985 845 75031 891
rect 75109 845 75155 891
rect 75233 845 75279 891
rect 75357 845 75403 891
rect 75481 845 75527 891
rect 75605 845 75651 891
rect 75729 845 75775 891
rect 75853 845 75899 891
rect 75977 845 76023 891
rect 76101 845 76147 891
rect 76225 845 76271 891
rect 76349 845 76395 891
rect 76473 845 76519 891
rect 76597 845 76643 891
rect 76721 845 76767 891
rect 76845 845 76891 891
rect 76969 845 77015 891
rect 77093 845 77139 891
rect 77217 845 77263 891
rect 77341 845 77387 891
rect 77465 845 77511 891
rect 77589 845 77635 891
rect 77713 845 77759 891
rect 77837 845 77883 891
rect 77961 845 78007 891
rect 78085 845 78131 891
rect 78209 845 78255 891
rect 78333 845 78379 891
rect 78457 845 78503 891
rect 78581 845 78627 891
rect 78705 845 78751 891
rect 78829 845 78875 891
rect 78953 845 78999 891
rect 79077 845 79123 891
rect 79201 845 79247 891
rect 79325 845 79371 891
rect 79449 845 79495 891
rect 79573 845 79619 891
rect 79697 845 79743 891
rect 79821 845 79867 891
rect 79945 845 79991 891
rect 80069 845 80115 891
rect 80193 845 80239 891
rect 80317 845 80363 891
rect 80441 845 80487 891
rect 80565 845 80611 891
rect 80689 845 80735 891
rect 80813 845 80859 891
rect 80937 845 80983 891
rect 81061 845 81107 891
rect 81185 845 81231 891
rect 81309 845 81355 891
rect 81433 845 81479 891
rect 81557 845 81603 891
rect 81681 845 81727 891
rect 81805 845 81851 891
rect 81929 845 81975 891
rect 82053 845 82099 891
rect 82177 845 82223 891
rect 82301 845 82347 891
rect 82425 845 82471 891
rect 82549 845 82595 891
rect 82673 845 82719 891
rect 82797 845 82843 891
rect 82921 845 82967 891
rect 83045 845 83091 891
rect 83169 845 83215 891
rect 83293 845 83339 891
rect 83417 845 83463 891
rect 83541 845 83587 891
rect 83665 845 83711 891
rect 83789 845 83835 891
rect 83913 845 83959 891
rect 84037 845 84083 891
rect 84161 845 84207 891
rect 84285 845 84331 891
rect 84409 845 84455 891
rect 84533 845 84579 891
rect 84657 845 84703 891
rect 84781 845 84827 891
rect 84905 845 84951 891
rect 85029 845 85075 891
rect 85153 845 85199 891
rect 85277 845 85323 891
rect 85401 845 85447 891
rect 85525 845 85571 891
rect 85649 845 85695 891
rect 89 721 135 767
rect 213 721 259 767
rect 337 721 383 767
rect 461 721 507 767
rect 585 721 631 767
rect 709 721 755 767
rect 833 721 879 767
rect 957 721 1003 767
rect 1081 721 1127 767
rect 1205 721 1251 767
rect 1329 721 1375 767
rect 1453 721 1499 767
rect 1577 721 1623 767
rect 1701 721 1747 767
rect 1825 721 1871 767
rect 1949 721 1995 767
rect 2073 721 2119 767
rect 2197 721 2243 767
rect 2321 721 2367 767
rect 2445 721 2491 767
rect 2569 721 2615 767
rect 2693 721 2739 767
rect 2817 721 2863 767
rect 2941 721 2987 767
rect 3065 721 3111 767
rect 3189 721 3235 767
rect 3313 721 3359 767
rect 3437 721 3483 767
rect 3561 721 3607 767
rect 3685 721 3731 767
rect 3809 721 3855 767
rect 3933 721 3979 767
rect 4057 721 4103 767
rect 4181 721 4227 767
rect 4305 721 4351 767
rect 4429 721 4475 767
rect 4553 721 4599 767
rect 4677 721 4723 767
rect 4801 721 4847 767
rect 4925 721 4971 767
rect 5049 721 5095 767
rect 5173 721 5219 767
rect 5297 721 5343 767
rect 5421 721 5467 767
rect 5545 721 5591 767
rect 5669 721 5715 767
rect 5793 721 5839 767
rect 5917 721 5963 767
rect 6041 721 6087 767
rect 6165 721 6211 767
rect 6289 721 6335 767
rect 6413 721 6459 767
rect 6537 721 6583 767
rect 6661 721 6707 767
rect 6785 721 6831 767
rect 6909 721 6955 767
rect 7033 721 7079 767
rect 7157 721 7203 767
rect 7281 721 7327 767
rect 7405 721 7451 767
rect 7529 721 7575 767
rect 7653 721 7699 767
rect 7777 721 7823 767
rect 7901 721 7947 767
rect 8025 721 8071 767
rect 8149 721 8195 767
rect 8273 721 8319 767
rect 8397 721 8443 767
rect 8521 721 8567 767
rect 8645 721 8691 767
rect 8769 721 8815 767
rect 8893 721 8939 767
rect 9017 721 9063 767
rect 9141 721 9187 767
rect 9265 721 9311 767
rect 9389 721 9435 767
rect 9513 721 9559 767
rect 9637 721 9683 767
rect 9761 721 9807 767
rect 9885 721 9931 767
rect 10009 721 10055 767
rect 10133 721 10179 767
rect 10257 721 10303 767
rect 10381 721 10427 767
rect 10505 721 10551 767
rect 10629 721 10675 767
rect 10753 721 10799 767
rect 10877 721 10923 767
rect 11001 721 11047 767
rect 11125 721 11171 767
rect 11249 721 11295 767
rect 11373 721 11419 767
rect 11497 721 11543 767
rect 11621 721 11667 767
rect 11745 721 11791 767
rect 11869 721 11915 767
rect 11993 721 12039 767
rect 12117 721 12163 767
rect 12241 721 12287 767
rect 12365 721 12411 767
rect 12489 721 12535 767
rect 12613 721 12659 767
rect 12737 721 12783 767
rect 12861 721 12907 767
rect 12985 721 13031 767
rect 13109 721 13155 767
rect 13233 721 13279 767
rect 13357 721 13403 767
rect 13481 721 13527 767
rect 13605 721 13651 767
rect 13729 721 13775 767
rect 13853 721 13899 767
rect 13977 721 14023 767
rect 14101 721 14147 767
rect 14225 721 14271 767
rect 14349 721 14395 767
rect 14473 721 14519 767
rect 14597 721 14643 767
rect 14721 721 14767 767
rect 14845 721 14891 767
rect 14969 721 15015 767
rect 15093 721 15139 767
rect 15217 721 15263 767
rect 15341 721 15387 767
rect 15465 721 15511 767
rect 15589 721 15635 767
rect 15713 721 15759 767
rect 15837 721 15883 767
rect 15961 721 16007 767
rect 16085 721 16131 767
rect 16209 721 16255 767
rect 16333 721 16379 767
rect 16457 721 16503 767
rect 16581 721 16627 767
rect 16705 721 16751 767
rect 16829 721 16875 767
rect 16953 721 16999 767
rect 17077 721 17123 767
rect 17201 721 17247 767
rect 17325 721 17371 767
rect 17449 721 17495 767
rect 17573 721 17619 767
rect 17697 721 17743 767
rect 17821 721 17867 767
rect 17945 721 17991 767
rect 18069 721 18115 767
rect 18193 721 18239 767
rect 18317 721 18363 767
rect 18441 721 18487 767
rect 18565 721 18611 767
rect 18689 721 18735 767
rect 18813 721 18859 767
rect 18937 721 18983 767
rect 19061 721 19107 767
rect 19185 721 19231 767
rect 19309 721 19355 767
rect 19433 721 19479 767
rect 19557 721 19603 767
rect 19681 721 19727 767
rect 19805 721 19851 767
rect 19929 721 19975 767
rect 20053 721 20099 767
rect 20177 721 20223 767
rect 20301 721 20347 767
rect 20425 721 20471 767
rect 20549 721 20595 767
rect 20673 721 20719 767
rect 20797 721 20843 767
rect 20921 721 20967 767
rect 21045 721 21091 767
rect 21169 721 21215 767
rect 21293 721 21339 767
rect 21417 721 21463 767
rect 21541 721 21587 767
rect 21665 721 21711 767
rect 21789 721 21835 767
rect 21913 721 21959 767
rect 22037 721 22083 767
rect 22161 721 22207 767
rect 22285 721 22331 767
rect 22409 721 22455 767
rect 22533 721 22579 767
rect 22657 721 22703 767
rect 22781 721 22827 767
rect 22905 721 22951 767
rect 23029 721 23075 767
rect 23153 721 23199 767
rect 23277 721 23323 767
rect 23401 721 23447 767
rect 23525 721 23571 767
rect 23649 721 23695 767
rect 23773 721 23819 767
rect 23897 721 23943 767
rect 24021 721 24067 767
rect 24145 721 24191 767
rect 24269 721 24315 767
rect 24393 721 24439 767
rect 24517 721 24563 767
rect 24641 721 24687 767
rect 24765 721 24811 767
rect 24889 721 24935 767
rect 25013 721 25059 767
rect 25137 721 25183 767
rect 25261 721 25307 767
rect 25385 721 25431 767
rect 25509 721 25555 767
rect 25633 721 25679 767
rect 25757 721 25803 767
rect 25881 721 25927 767
rect 26005 721 26051 767
rect 26129 721 26175 767
rect 26253 721 26299 767
rect 26377 721 26423 767
rect 26501 721 26547 767
rect 26625 721 26671 767
rect 26749 721 26795 767
rect 26873 721 26919 767
rect 26997 721 27043 767
rect 27121 721 27167 767
rect 27245 721 27291 767
rect 27369 721 27415 767
rect 27493 721 27539 767
rect 27617 721 27663 767
rect 27741 721 27787 767
rect 27865 721 27911 767
rect 27989 721 28035 767
rect 28113 721 28159 767
rect 28237 721 28283 767
rect 28361 721 28407 767
rect 28485 721 28531 767
rect 28609 721 28655 767
rect 28733 721 28779 767
rect 28857 721 28903 767
rect 28981 721 29027 767
rect 29105 721 29151 767
rect 29229 721 29275 767
rect 29353 721 29399 767
rect 29477 721 29523 767
rect 29601 721 29647 767
rect 29725 721 29771 767
rect 29849 721 29895 767
rect 29973 721 30019 767
rect 30097 721 30143 767
rect 30221 721 30267 767
rect 30345 721 30391 767
rect 30469 721 30515 767
rect 30593 721 30639 767
rect 30717 721 30763 767
rect 30841 721 30887 767
rect 30965 721 31011 767
rect 31089 721 31135 767
rect 31213 721 31259 767
rect 31337 721 31383 767
rect 31461 721 31507 767
rect 31585 721 31631 767
rect 31709 721 31755 767
rect 31833 721 31879 767
rect 31957 721 32003 767
rect 32081 721 32127 767
rect 32205 721 32251 767
rect 32329 721 32375 767
rect 32453 721 32499 767
rect 32577 721 32623 767
rect 32701 721 32747 767
rect 32825 721 32871 767
rect 32949 721 32995 767
rect 33073 721 33119 767
rect 33197 721 33243 767
rect 33321 721 33367 767
rect 33445 721 33491 767
rect 33569 721 33615 767
rect 33693 721 33739 767
rect 33817 721 33863 767
rect 33941 721 33987 767
rect 34065 721 34111 767
rect 34189 721 34235 767
rect 34313 721 34359 767
rect 34437 721 34483 767
rect 34561 721 34607 767
rect 34685 721 34731 767
rect 34809 721 34855 767
rect 34933 721 34979 767
rect 35057 721 35103 767
rect 35181 721 35227 767
rect 35305 721 35351 767
rect 35429 721 35475 767
rect 35553 721 35599 767
rect 35677 721 35723 767
rect 35801 721 35847 767
rect 35925 721 35971 767
rect 36049 721 36095 767
rect 36173 721 36219 767
rect 36297 721 36343 767
rect 36421 721 36467 767
rect 36545 721 36591 767
rect 36669 721 36715 767
rect 36793 721 36839 767
rect 36917 721 36963 767
rect 37041 721 37087 767
rect 37165 721 37211 767
rect 37289 721 37335 767
rect 37413 721 37459 767
rect 37537 721 37583 767
rect 37661 721 37707 767
rect 37785 721 37831 767
rect 37909 721 37955 767
rect 38033 721 38079 767
rect 38157 721 38203 767
rect 38281 721 38327 767
rect 38405 721 38451 767
rect 38529 721 38575 767
rect 38653 721 38699 767
rect 38777 721 38823 767
rect 38901 721 38947 767
rect 39025 721 39071 767
rect 39149 721 39195 767
rect 39273 721 39319 767
rect 39397 721 39443 767
rect 39521 721 39567 767
rect 39645 721 39691 767
rect 39769 721 39815 767
rect 39893 721 39939 767
rect 40017 721 40063 767
rect 40141 721 40187 767
rect 40265 721 40311 767
rect 40389 721 40435 767
rect 40513 721 40559 767
rect 40637 721 40683 767
rect 40761 721 40807 767
rect 40885 721 40931 767
rect 41009 721 41055 767
rect 41133 721 41179 767
rect 41257 721 41303 767
rect 41381 721 41427 767
rect 41505 721 41551 767
rect 41629 721 41675 767
rect 41753 721 41799 767
rect 41877 721 41923 767
rect 42001 721 42047 767
rect 42125 721 42171 767
rect 42249 721 42295 767
rect 42373 721 42419 767
rect 42497 721 42543 767
rect 42621 721 42667 767
rect 42745 721 42791 767
rect 42869 721 42915 767
rect 42993 721 43039 767
rect 43117 721 43163 767
rect 43241 721 43287 767
rect 43365 721 43411 767
rect 43489 721 43535 767
rect 43613 721 43659 767
rect 43737 721 43783 767
rect 43861 721 43907 767
rect 43985 721 44031 767
rect 44109 721 44155 767
rect 44233 721 44279 767
rect 44357 721 44403 767
rect 44481 721 44527 767
rect 44605 721 44651 767
rect 44729 721 44775 767
rect 44853 721 44899 767
rect 44977 721 45023 767
rect 45101 721 45147 767
rect 45225 721 45271 767
rect 45349 721 45395 767
rect 45473 721 45519 767
rect 45597 721 45643 767
rect 45721 721 45767 767
rect 45845 721 45891 767
rect 45969 721 46015 767
rect 46093 721 46139 767
rect 46217 721 46263 767
rect 46341 721 46387 767
rect 46465 721 46511 767
rect 46589 721 46635 767
rect 46713 721 46759 767
rect 46837 721 46883 767
rect 46961 721 47007 767
rect 47085 721 47131 767
rect 47209 721 47255 767
rect 47333 721 47379 767
rect 47457 721 47503 767
rect 47581 721 47627 767
rect 47705 721 47751 767
rect 47829 721 47875 767
rect 47953 721 47999 767
rect 48077 721 48123 767
rect 48201 721 48247 767
rect 48325 721 48371 767
rect 48449 721 48495 767
rect 48573 721 48619 767
rect 48697 721 48743 767
rect 48821 721 48867 767
rect 48945 721 48991 767
rect 49069 721 49115 767
rect 49193 721 49239 767
rect 49317 721 49363 767
rect 49441 721 49487 767
rect 49565 721 49611 767
rect 49689 721 49735 767
rect 49813 721 49859 767
rect 49937 721 49983 767
rect 50061 721 50107 767
rect 50185 721 50231 767
rect 50309 721 50355 767
rect 50433 721 50479 767
rect 50557 721 50603 767
rect 50681 721 50727 767
rect 50805 721 50851 767
rect 50929 721 50975 767
rect 51053 721 51099 767
rect 51177 721 51223 767
rect 51301 721 51347 767
rect 51425 721 51471 767
rect 51549 721 51595 767
rect 51673 721 51719 767
rect 51797 721 51843 767
rect 51921 721 51967 767
rect 52045 721 52091 767
rect 52169 721 52215 767
rect 52293 721 52339 767
rect 52417 721 52463 767
rect 52541 721 52587 767
rect 52665 721 52711 767
rect 52789 721 52835 767
rect 52913 721 52959 767
rect 53037 721 53083 767
rect 53161 721 53207 767
rect 53285 721 53331 767
rect 53409 721 53455 767
rect 53533 721 53579 767
rect 53657 721 53703 767
rect 53781 721 53827 767
rect 53905 721 53951 767
rect 54029 721 54075 767
rect 54153 721 54199 767
rect 54277 721 54323 767
rect 54401 721 54447 767
rect 54525 721 54571 767
rect 54649 721 54695 767
rect 54773 721 54819 767
rect 54897 721 54943 767
rect 55021 721 55067 767
rect 55145 721 55191 767
rect 55269 721 55315 767
rect 55393 721 55439 767
rect 55517 721 55563 767
rect 55641 721 55687 767
rect 55765 721 55811 767
rect 55889 721 55935 767
rect 56013 721 56059 767
rect 56137 721 56183 767
rect 56261 721 56307 767
rect 56385 721 56431 767
rect 56509 721 56555 767
rect 56633 721 56679 767
rect 56757 721 56803 767
rect 56881 721 56927 767
rect 57005 721 57051 767
rect 57129 721 57175 767
rect 57253 721 57299 767
rect 57377 721 57423 767
rect 57501 721 57547 767
rect 57625 721 57671 767
rect 57749 721 57795 767
rect 57873 721 57919 767
rect 57997 721 58043 767
rect 58121 721 58167 767
rect 58245 721 58291 767
rect 58369 721 58415 767
rect 58493 721 58539 767
rect 58617 721 58663 767
rect 58741 721 58787 767
rect 58865 721 58911 767
rect 58989 721 59035 767
rect 59113 721 59159 767
rect 59237 721 59283 767
rect 59361 721 59407 767
rect 59485 721 59531 767
rect 59609 721 59655 767
rect 59733 721 59779 767
rect 59857 721 59903 767
rect 59981 721 60027 767
rect 60105 721 60151 767
rect 60229 721 60275 767
rect 60353 721 60399 767
rect 60477 721 60523 767
rect 60601 721 60647 767
rect 60725 721 60771 767
rect 60849 721 60895 767
rect 60973 721 61019 767
rect 61097 721 61143 767
rect 61221 721 61267 767
rect 61345 721 61391 767
rect 61469 721 61515 767
rect 61593 721 61639 767
rect 61717 721 61763 767
rect 61841 721 61887 767
rect 61965 721 62011 767
rect 62089 721 62135 767
rect 62213 721 62259 767
rect 62337 721 62383 767
rect 62461 721 62507 767
rect 62585 721 62631 767
rect 62709 721 62755 767
rect 62833 721 62879 767
rect 62957 721 63003 767
rect 63081 721 63127 767
rect 63205 721 63251 767
rect 63329 721 63375 767
rect 63453 721 63499 767
rect 63577 721 63623 767
rect 63701 721 63747 767
rect 63825 721 63871 767
rect 63949 721 63995 767
rect 64073 721 64119 767
rect 64197 721 64243 767
rect 64321 721 64367 767
rect 64445 721 64491 767
rect 64569 721 64615 767
rect 64693 721 64739 767
rect 64817 721 64863 767
rect 64941 721 64987 767
rect 65065 721 65111 767
rect 65189 721 65235 767
rect 65313 721 65359 767
rect 65437 721 65483 767
rect 65561 721 65607 767
rect 65685 721 65731 767
rect 65809 721 65855 767
rect 65933 721 65979 767
rect 66057 721 66103 767
rect 66181 721 66227 767
rect 66305 721 66351 767
rect 66429 721 66475 767
rect 66553 721 66599 767
rect 66677 721 66723 767
rect 66801 721 66847 767
rect 66925 721 66971 767
rect 67049 721 67095 767
rect 67173 721 67219 767
rect 67297 721 67343 767
rect 67421 721 67467 767
rect 67545 721 67591 767
rect 67669 721 67715 767
rect 67793 721 67839 767
rect 67917 721 67963 767
rect 68041 721 68087 767
rect 68165 721 68211 767
rect 68289 721 68335 767
rect 68413 721 68459 767
rect 68537 721 68583 767
rect 68661 721 68707 767
rect 68785 721 68831 767
rect 68909 721 68955 767
rect 69033 721 69079 767
rect 69157 721 69203 767
rect 69281 721 69327 767
rect 69405 721 69451 767
rect 69529 721 69575 767
rect 69653 721 69699 767
rect 69777 721 69823 767
rect 69901 721 69947 767
rect 70025 721 70071 767
rect 70149 721 70195 767
rect 70273 721 70319 767
rect 70397 721 70443 767
rect 70521 721 70567 767
rect 70645 721 70691 767
rect 70769 721 70815 767
rect 70893 721 70939 767
rect 71017 721 71063 767
rect 71141 721 71187 767
rect 71265 721 71311 767
rect 71389 721 71435 767
rect 71513 721 71559 767
rect 71637 721 71683 767
rect 71761 721 71807 767
rect 71885 721 71931 767
rect 72009 721 72055 767
rect 72133 721 72179 767
rect 72257 721 72303 767
rect 72381 721 72427 767
rect 72505 721 72551 767
rect 72629 721 72675 767
rect 72753 721 72799 767
rect 72877 721 72923 767
rect 73001 721 73047 767
rect 73125 721 73171 767
rect 73249 721 73295 767
rect 73373 721 73419 767
rect 73497 721 73543 767
rect 73621 721 73667 767
rect 73745 721 73791 767
rect 73869 721 73915 767
rect 73993 721 74039 767
rect 74117 721 74163 767
rect 74241 721 74287 767
rect 74365 721 74411 767
rect 74489 721 74535 767
rect 74613 721 74659 767
rect 74737 721 74783 767
rect 74861 721 74907 767
rect 74985 721 75031 767
rect 75109 721 75155 767
rect 75233 721 75279 767
rect 75357 721 75403 767
rect 75481 721 75527 767
rect 75605 721 75651 767
rect 75729 721 75775 767
rect 75853 721 75899 767
rect 75977 721 76023 767
rect 76101 721 76147 767
rect 76225 721 76271 767
rect 76349 721 76395 767
rect 76473 721 76519 767
rect 76597 721 76643 767
rect 76721 721 76767 767
rect 76845 721 76891 767
rect 76969 721 77015 767
rect 77093 721 77139 767
rect 77217 721 77263 767
rect 77341 721 77387 767
rect 77465 721 77511 767
rect 77589 721 77635 767
rect 77713 721 77759 767
rect 77837 721 77883 767
rect 77961 721 78007 767
rect 78085 721 78131 767
rect 78209 721 78255 767
rect 78333 721 78379 767
rect 78457 721 78503 767
rect 78581 721 78627 767
rect 78705 721 78751 767
rect 78829 721 78875 767
rect 78953 721 78999 767
rect 79077 721 79123 767
rect 79201 721 79247 767
rect 79325 721 79371 767
rect 79449 721 79495 767
rect 79573 721 79619 767
rect 79697 721 79743 767
rect 79821 721 79867 767
rect 79945 721 79991 767
rect 80069 721 80115 767
rect 80193 721 80239 767
rect 80317 721 80363 767
rect 80441 721 80487 767
rect 80565 721 80611 767
rect 80689 721 80735 767
rect 80813 721 80859 767
rect 80937 721 80983 767
rect 81061 721 81107 767
rect 81185 721 81231 767
rect 81309 721 81355 767
rect 81433 721 81479 767
rect 81557 721 81603 767
rect 81681 721 81727 767
rect 81805 721 81851 767
rect 81929 721 81975 767
rect 82053 721 82099 767
rect 82177 721 82223 767
rect 82301 721 82347 767
rect 82425 721 82471 767
rect 82549 721 82595 767
rect 82673 721 82719 767
rect 82797 721 82843 767
rect 82921 721 82967 767
rect 83045 721 83091 767
rect 83169 721 83215 767
rect 83293 721 83339 767
rect 83417 721 83463 767
rect 83541 721 83587 767
rect 83665 721 83711 767
rect 83789 721 83835 767
rect 83913 721 83959 767
rect 84037 721 84083 767
rect 84161 721 84207 767
rect 84285 721 84331 767
rect 84409 721 84455 767
rect 84533 721 84579 767
rect 84657 721 84703 767
rect 84781 721 84827 767
rect 84905 721 84951 767
rect 85029 721 85075 767
rect 85153 721 85199 767
rect 85277 721 85323 767
rect 85401 721 85447 767
rect 85525 721 85571 767
rect 85649 721 85695 767
rect 89 597 135 643
rect 213 597 259 643
rect 337 597 383 643
rect 461 597 507 643
rect 585 597 631 643
rect 709 597 755 643
rect 833 597 879 643
rect 957 597 1003 643
rect 1081 597 1127 643
rect 1205 597 1251 643
rect 1329 597 1375 643
rect 1453 597 1499 643
rect 1577 597 1623 643
rect 1701 597 1747 643
rect 1825 597 1871 643
rect 1949 597 1995 643
rect 2073 597 2119 643
rect 2197 597 2243 643
rect 2321 597 2367 643
rect 2445 597 2491 643
rect 2569 597 2615 643
rect 2693 597 2739 643
rect 2817 597 2863 643
rect 2941 597 2987 643
rect 3065 597 3111 643
rect 3189 597 3235 643
rect 3313 597 3359 643
rect 3437 597 3483 643
rect 3561 597 3607 643
rect 3685 597 3731 643
rect 3809 597 3855 643
rect 3933 597 3979 643
rect 4057 597 4103 643
rect 4181 597 4227 643
rect 4305 597 4351 643
rect 4429 597 4475 643
rect 4553 597 4599 643
rect 4677 597 4723 643
rect 4801 597 4847 643
rect 4925 597 4971 643
rect 5049 597 5095 643
rect 5173 597 5219 643
rect 5297 597 5343 643
rect 5421 597 5467 643
rect 5545 597 5591 643
rect 5669 597 5715 643
rect 5793 597 5839 643
rect 5917 597 5963 643
rect 6041 597 6087 643
rect 6165 597 6211 643
rect 6289 597 6335 643
rect 6413 597 6459 643
rect 6537 597 6583 643
rect 6661 597 6707 643
rect 6785 597 6831 643
rect 6909 597 6955 643
rect 7033 597 7079 643
rect 7157 597 7203 643
rect 7281 597 7327 643
rect 7405 597 7451 643
rect 7529 597 7575 643
rect 7653 597 7699 643
rect 7777 597 7823 643
rect 7901 597 7947 643
rect 8025 597 8071 643
rect 8149 597 8195 643
rect 8273 597 8319 643
rect 8397 597 8443 643
rect 8521 597 8567 643
rect 8645 597 8691 643
rect 8769 597 8815 643
rect 8893 597 8939 643
rect 9017 597 9063 643
rect 9141 597 9187 643
rect 9265 597 9311 643
rect 9389 597 9435 643
rect 9513 597 9559 643
rect 9637 597 9683 643
rect 9761 597 9807 643
rect 9885 597 9931 643
rect 10009 597 10055 643
rect 10133 597 10179 643
rect 10257 597 10303 643
rect 10381 597 10427 643
rect 10505 597 10551 643
rect 10629 597 10675 643
rect 10753 597 10799 643
rect 10877 597 10923 643
rect 11001 597 11047 643
rect 11125 597 11171 643
rect 11249 597 11295 643
rect 11373 597 11419 643
rect 11497 597 11543 643
rect 11621 597 11667 643
rect 11745 597 11791 643
rect 11869 597 11915 643
rect 11993 597 12039 643
rect 12117 597 12163 643
rect 12241 597 12287 643
rect 12365 597 12411 643
rect 12489 597 12535 643
rect 12613 597 12659 643
rect 12737 597 12783 643
rect 12861 597 12907 643
rect 12985 597 13031 643
rect 13109 597 13155 643
rect 13233 597 13279 643
rect 13357 597 13403 643
rect 13481 597 13527 643
rect 13605 597 13651 643
rect 13729 597 13775 643
rect 13853 597 13899 643
rect 13977 597 14023 643
rect 14101 597 14147 643
rect 14225 597 14271 643
rect 14349 597 14395 643
rect 14473 597 14519 643
rect 14597 597 14643 643
rect 14721 597 14767 643
rect 14845 597 14891 643
rect 14969 597 15015 643
rect 15093 597 15139 643
rect 15217 597 15263 643
rect 15341 597 15387 643
rect 15465 597 15511 643
rect 15589 597 15635 643
rect 15713 597 15759 643
rect 15837 597 15883 643
rect 15961 597 16007 643
rect 16085 597 16131 643
rect 16209 597 16255 643
rect 16333 597 16379 643
rect 16457 597 16503 643
rect 16581 597 16627 643
rect 16705 597 16751 643
rect 16829 597 16875 643
rect 16953 597 16999 643
rect 17077 597 17123 643
rect 17201 597 17247 643
rect 17325 597 17371 643
rect 17449 597 17495 643
rect 17573 597 17619 643
rect 17697 597 17743 643
rect 17821 597 17867 643
rect 17945 597 17991 643
rect 18069 597 18115 643
rect 18193 597 18239 643
rect 18317 597 18363 643
rect 18441 597 18487 643
rect 18565 597 18611 643
rect 18689 597 18735 643
rect 18813 597 18859 643
rect 18937 597 18983 643
rect 19061 597 19107 643
rect 19185 597 19231 643
rect 19309 597 19355 643
rect 19433 597 19479 643
rect 19557 597 19603 643
rect 19681 597 19727 643
rect 19805 597 19851 643
rect 19929 597 19975 643
rect 20053 597 20099 643
rect 20177 597 20223 643
rect 20301 597 20347 643
rect 20425 597 20471 643
rect 20549 597 20595 643
rect 20673 597 20719 643
rect 20797 597 20843 643
rect 20921 597 20967 643
rect 21045 597 21091 643
rect 21169 597 21215 643
rect 21293 597 21339 643
rect 21417 597 21463 643
rect 21541 597 21587 643
rect 21665 597 21711 643
rect 21789 597 21835 643
rect 21913 597 21959 643
rect 22037 597 22083 643
rect 22161 597 22207 643
rect 22285 597 22331 643
rect 22409 597 22455 643
rect 22533 597 22579 643
rect 22657 597 22703 643
rect 22781 597 22827 643
rect 22905 597 22951 643
rect 23029 597 23075 643
rect 23153 597 23199 643
rect 23277 597 23323 643
rect 23401 597 23447 643
rect 23525 597 23571 643
rect 23649 597 23695 643
rect 23773 597 23819 643
rect 23897 597 23943 643
rect 24021 597 24067 643
rect 24145 597 24191 643
rect 24269 597 24315 643
rect 24393 597 24439 643
rect 24517 597 24563 643
rect 24641 597 24687 643
rect 24765 597 24811 643
rect 24889 597 24935 643
rect 25013 597 25059 643
rect 25137 597 25183 643
rect 25261 597 25307 643
rect 25385 597 25431 643
rect 25509 597 25555 643
rect 25633 597 25679 643
rect 25757 597 25803 643
rect 25881 597 25927 643
rect 26005 597 26051 643
rect 26129 597 26175 643
rect 26253 597 26299 643
rect 26377 597 26423 643
rect 26501 597 26547 643
rect 26625 597 26671 643
rect 26749 597 26795 643
rect 26873 597 26919 643
rect 26997 597 27043 643
rect 27121 597 27167 643
rect 27245 597 27291 643
rect 27369 597 27415 643
rect 27493 597 27539 643
rect 27617 597 27663 643
rect 27741 597 27787 643
rect 27865 597 27911 643
rect 27989 597 28035 643
rect 28113 597 28159 643
rect 28237 597 28283 643
rect 28361 597 28407 643
rect 28485 597 28531 643
rect 28609 597 28655 643
rect 28733 597 28779 643
rect 28857 597 28903 643
rect 28981 597 29027 643
rect 29105 597 29151 643
rect 29229 597 29275 643
rect 29353 597 29399 643
rect 29477 597 29523 643
rect 29601 597 29647 643
rect 29725 597 29771 643
rect 29849 597 29895 643
rect 29973 597 30019 643
rect 30097 597 30143 643
rect 30221 597 30267 643
rect 30345 597 30391 643
rect 30469 597 30515 643
rect 30593 597 30639 643
rect 30717 597 30763 643
rect 30841 597 30887 643
rect 30965 597 31011 643
rect 31089 597 31135 643
rect 31213 597 31259 643
rect 31337 597 31383 643
rect 31461 597 31507 643
rect 31585 597 31631 643
rect 31709 597 31755 643
rect 31833 597 31879 643
rect 31957 597 32003 643
rect 32081 597 32127 643
rect 32205 597 32251 643
rect 32329 597 32375 643
rect 32453 597 32499 643
rect 32577 597 32623 643
rect 32701 597 32747 643
rect 32825 597 32871 643
rect 32949 597 32995 643
rect 33073 597 33119 643
rect 33197 597 33243 643
rect 33321 597 33367 643
rect 33445 597 33491 643
rect 33569 597 33615 643
rect 33693 597 33739 643
rect 33817 597 33863 643
rect 33941 597 33987 643
rect 34065 597 34111 643
rect 34189 597 34235 643
rect 34313 597 34359 643
rect 34437 597 34483 643
rect 34561 597 34607 643
rect 34685 597 34731 643
rect 34809 597 34855 643
rect 34933 597 34979 643
rect 35057 597 35103 643
rect 35181 597 35227 643
rect 35305 597 35351 643
rect 35429 597 35475 643
rect 35553 597 35599 643
rect 35677 597 35723 643
rect 35801 597 35847 643
rect 35925 597 35971 643
rect 36049 597 36095 643
rect 36173 597 36219 643
rect 36297 597 36343 643
rect 36421 597 36467 643
rect 36545 597 36591 643
rect 36669 597 36715 643
rect 36793 597 36839 643
rect 36917 597 36963 643
rect 37041 597 37087 643
rect 37165 597 37211 643
rect 37289 597 37335 643
rect 37413 597 37459 643
rect 37537 597 37583 643
rect 37661 597 37707 643
rect 37785 597 37831 643
rect 37909 597 37955 643
rect 38033 597 38079 643
rect 38157 597 38203 643
rect 38281 597 38327 643
rect 38405 597 38451 643
rect 38529 597 38575 643
rect 38653 597 38699 643
rect 38777 597 38823 643
rect 38901 597 38947 643
rect 39025 597 39071 643
rect 39149 597 39195 643
rect 39273 597 39319 643
rect 39397 597 39443 643
rect 39521 597 39567 643
rect 39645 597 39691 643
rect 39769 597 39815 643
rect 39893 597 39939 643
rect 40017 597 40063 643
rect 40141 597 40187 643
rect 40265 597 40311 643
rect 40389 597 40435 643
rect 40513 597 40559 643
rect 40637 597 40683 643
rect 40761 597 40807 643
rect 40885 597 40931 643
rect 41009 597 41055 643
rect 41133 597 41179 643
rect 41257 597 41303 643
rect 41381 597 41427 643
rect 41505 597 41551 643
rect 41629 597 41675 643
rect 41753 597 41799 643
rect 41877 597 41923 643
rect 42001 597 42047 643
rect 42125 597 42171 643
rect 42249 597 42295 643
rect 42373 597 42419 643
rect 42497 597 42543 643
rect 42621 597 42667 643
rect 42745 597 42791 643
rect 42869 597 42915 643
rect 42993 597 43039 643
rect 43117 597 43163 643
rect 43241 597 43287 643
rect 43365 597 43411 643
rect 43489 597 43535 643
rect 43613 597 43659 643
rect 43737 597 43783 643
rect 43861 597 43907 643
rect 43985 597 44031 643
rect 44109 597 44155 643
rect 44233 597 44279 643
rect 44357 597 44403 643
rect 44481 597 44527 643
rect 44605 597 44651 643
rect 44729 597 44775 643
rect 44853 597 44899 643
rect 44977 597 45023 643
rect 45101 597 45147 643
rect 45225 597 45271 643
rect 45349 597 45395 643
rect 45473 597 45519 643
rect 45597 597 45643 643
rect 45721 597 45767 643
rect 45845 597 45891 643
rect 45969 597 46015 643
rect 46093 597 46139 643
rect 46217 597 46263 643
rect 46341 597 46387 643
rect 46465 597 46511 643
rect 46589 597 46635 643
rect 46713 597 46759 643
rect 46837 597 46883 643
rect 46961 597 47007 643
rect 47085 597 47131 643
rect 47209 597 47255 643
rect 47333 597 47379 643
rect 47457 597 47503 643
rect 47581 597 47627 643
rect 47705 597 47751 643
rect 47829 597 47875 643
rect 47953 597 47999 643
rect 48077 597 48123 643
rect 48201 597 48247 643
rect 48325 597 48371 643
rect 48449 597 48495 643
rect 48573 597 48619 643
rect 48697 597 48743 643
rect 48821 597 48867 643
rect 48945 597 48991 643
rect 49069 597 49115 643
rect 49193 597 49239 643
rect 49317 597 49363 643
rect 49441 597 49487 643
rect 49565 597 49611 643
rect 49689 597 49735 643
rect 49813 597 49859 643
rect 49937 597 49983 643
rect 50061 597 50107 643
rect 50185 597 50231 643
rect 50309 597 50355 643
rect 50433 597 50479 643
rect 50557 597 50603 643
rect 50681 597 50727 643
rect 50805 597 50851 643
rect 50929 597 50975 643
rect 51053 597 51099 643
rect 51177 597 51223 643
rect 51301 597 51347 643
rect 51425 597 51471 643
rect 51549 597 51595 643
rect 51673 597 51719 643
rect 51797 597 51843 643
rect 51921 597 51967 643
rect 52045 597 52091 643
rect 52169 597 52215 643
rect 52293 597 52339 643
rect 52417 597 52463 643
rect 52541 597 52587 643
rect 52665 597 52711 643
rect 52789 597 52835 643
rect 52913 597 52959 643
rect 53037 597 53083 643
rect 53161 597 53207 643
rect 53285 597 53331 643
rect 53409 597 53455 643
rect 53533 597 53579 643
rect 53657 597 53703 643
rect 53781 597 53827 643
rect 53905 597 53951 643
rect 54029 597 54075 643
rect 54153 597 54199 643
rect 54277 597 54323 643
rect 54401 597 54447 643
rect 54525 597 54571 643
rect 54649 597 54695 643
rect 54773 597 54819 643
rect 54897 597 54943 643
rect 55021 597 55067 643
rect 55145 597 55191 643
rect 55269 597 55315 643
rect 55393 597 55439 643
rect 55517 597 55563 643
rect 55641 597 55687 643
rect 55765 597 55811 643
rect 55889 597 55935 643
rect 56013 597 56059 643
rect 56137 597 56183 643
rect 56261 597 56307 643
rect 56385 597 56431 643
rect 56509 597 56555 643
rect 56633 597 56679 643
rect 56757 597 56803 643
rect 56881 597 56927 643
rect 57005 597 57051 643
rect 57129 597 57175 643
rect 57253 597 57299 643
rect 57377 597 57423 643
rect 57501 597 57547 643
rect 57625 597 57671 643
rect 57749 597 57795 643
rect 57873 597 57919 643
rect 57997 597 58043 643
rect 58121 597 58167 643
rect 58245 597 58291 643
rect 58369 597 58415 643
rect 58493 597 58539 643
rect 58617 597 58663 643
rect 58741 597 58787 643
rect 58865 597 58911 643
rect 58989 597 59035 643
rect 59113 597 59159 643
rect 59237 597 59283 643
rect 59361 597 59407 643
rect 59485 597 59531 643
rect 59609 597 59655 643
rect 59733 597 59779 643
rect 59857 597 59903 643
rect 59981 597 60027 643
rect 60105 597 60151 643
rect 60229 597 60275 643
rect 60353 597 60399 643
rect 60477 597 60523 643
rect 60601 597 60647 643
rect 60725 597 60771 643
rect 60849 597 60895 643
rect 60973 597 61019 643
rect 61097 597 61143 643
rect 61221 597 61267 643
rect 61345 597 61391 643
rect 61469 597 61515 643
rect 61593 597 61639 643
rect 61717 597 61763 643
rect 61841 597 61887 643
rect 61965 597 62011 643
rect 62089 597 62135 643
rect 62213 597 62259 643
rect 62337 597 62383 643
rect 62461 597 62507 643
rect 62585 597 62631 643
rect 62709 597 62755 643
rect 62833 597 62879 643
rect 62957 597 63003 643
rect 63081 597 63127 643
rect 63205 597 63251 643
rect 63329 597 63375 643
rect 63453 597 63499 643
rect 63577 597 63623 643
rect 63701 597 63747 643
rect 63825 597 63871 643
rect 63949 597 63995 643
rect 64073 597 64119 643
rect 64197 597 64243 643
rect 64321 597 64367 643
rect 64445 597 64491 643
rect 64569 597 64615 643
rect 64693 597 64739 643
rect 64817 597 64863 643
rect 64941 597 64987 643
rect 65065 597 65111 643
rect 65189 597 65235 643
rect 65313 597 65359 643
rect 65437 597 65483 643
rect 65561 597 65607 643
rect 65685 597 65731 643
rect 65809 597 65855 643
rect 65933 597 65979 643
rect 66057 597 66103 643
rect 66181 597 66227 643
rect 66305 597 66351 643
rect 66429 597 66475 643
rect 66553 597 66599 643
rect 66677 597 66723 643
rect 66801 597 66847 643
rect 66925 597 66971 643
rect 67049 597 67095 643
rect 67173 597 67219 643
rect 67297 597 67343 643
rect 67421 597 67467 643
rect 67545 597 67591 643
rect 67669 597 67715 643
rect 67793 597 67839 643
rect 67917 597 67963 643
rect 68041 597 68087 643
rect 68165 597 68211 643
rect 68289 597 68335 643
rect 68413 597 68459 643
rect 68537 597 68583 643
rect 68661 597 68707 643
rect 68785 597 68831 643
rect 68909 597 68955 643
rect 69033 597 69079 643
rect 69157 597 69203 643
rect 69281 597 69327 643
rect 69405 597 69451 643
rect 69529 597 69575 643
rect 69653 597 69699 643
rect 69777 597 69823 643
rect 69901 597 69947 643
rect 70025 597 70071 643
rect 70149 597 70195 643
rect 70273 597 70319 643
rect 70397 597 70443 643
rect 70521 597 70567 643
rect 70645 597 70691 643
rect 70769 597 70815 643
rect 70893 597 70939 643
rect 71017 597 71063 643
rect 71141 597 71187 643
rect 71265 597 71311 643
rect 71389 597 71435 643
rect 71513 597 71559 643
rect 71637 597 71683 643
rect 71761 597 71807 643
rect 71885 597 71931 643
rect 72009 597 72055 643
rect 72133 597 72179 643
rect 72257 597 72303 643
rect 72381 597 72427 643
rect 72505 597 72551 643
rect 72629 597 72675 643
rect 72753 597 72799 643
rect 72877 597 72923 643
rect 73001 597 73047 643
rect 73125 597 73171 643
rect 73249 597 73295 643
rect 73373 597 73419 643
rect 73497 597 73543 643
rect 73621 597 73667 643
rect 73745 597 73791 643
rect 73869 597 73915 643
rect 73993 597 74039 643
rect 74117 597 74163 643
rect 74241 597 74287 643
rect 74365 597 74411 643
rect 74489 597 74535 643
rect 74613 597 74659 643
rect 74737 597 74783 643
rect 74861 597 74907 643
rect 74985 597 75031 643
rect 75109 597 75155 643
rect 75233 597 75279 643
rect 75357 597 75403 643
rect 75481 597 75527 643
rect 75605 597 75651 643
rect 75729 597 75775 643
rect 75853 597 75899 643
rect 75977 597 76023 643
rect 76101 597 76147 643
rect 76225 597 76271 643
rect 76349 597 76395 643
rect 76473 597 76519 643
rect 76597 597 76643 643
rect 76721 597 76767 643
rect 76845 597 76891 643
rect 76969 597 77015 643
rect 77093 597 77139 643
rect 77217 597 77263 643
rect 77341 597 77387 643
rect 77465 597 77511 643
rect 77589 597 77635 643
rect 77713 597 77759 643
rect 77837 597 77883 643
rect 77961 597 78007 643
rect 78085 597 78131 643
rect 78209 597 78255 643
rect 78333 597 78379 643
rect 78457 597 78503 643
rect 78581 597 78627 643
rect 78705 597 78751 643
rect 78829 597 78875 643
rect 78953 597 78999 643
rect 79077 597 79123 643
rect 79201 597 79247 643
rect 79325 597 79371 643
rect 79449 597 79495 643
rect 79573 597 79619 643
rect 79697 597 79743 643
rect 79821 597 79867 643
rect 79945 597 79991 643
rect 80069 597 80115 643
rect 80193 597 80239 643
rect 80317 597 80363 643
rect 80441 597 80487 643
rect 80565 597 80611 643
rect 80689 597 80735 643
rect 80813 597 80859 643
rect 80937 597 80983 643
rect 81061 597 81107 643
rect 81185 597 81231 643
rect 81309 597 81355 643
rect 81433 597 81479 643
rect 81557 597 81603 643
rect 81681 597 81727 643
rect 81805 597 81851 643
rect 81929 597 81975 643
rect 82053 597 82099 643
rect 82177 597 82223 643
rect 82301 597 82347 643
rect 82425 597 82471 643
rect 82549 597 82595 643
rect 82673 597 82719 643
rect 82797 597 82843 643
rect 82921 597 82967 643
rect 83045 597 83091 643
rect 83169 597 83215 643
rect 83293 597 83339 643
rect 83417 597 83463 643
rect 83541 597 83587 643
rect 83665 597 83711 643
rect 83789 597 83835 643
rect 83913 597 83959 643
rect 84037 597 84083 643
rect 84161 597 84207 643
rect 84285 597 84331 643
rect 84409 597 84455 643
rect 84533 597 84579 643
rect 84657 597 84703 643
rect 84781 597 84827 643
rect 84905 597 84951 643
rect 85029 597 85075 643
rect 85153 597 85199 643
rect 85277 597 85323 643
rect 85401 597 85447 643
rect 85525 597 85571 643
rect 85649 597 85695 643
<< metal1 >>
rect 0 53483 85706 53494
rect 0 53437 89 53483
rect 135 53437 213 53483
rect 259 53437 337 53483
rect 383 53437 461 53483
rect 507 53437 585 53483
rect 631 53437 709 53483
rect 755 53437 833 53483
rect 879 53437 957 53483
rect 1003 53437 1081 53483
rect 1127 53437 1205 53483
rect 1251 53437 1329 53483
rect 1375 53437 1453 53483
rect 1499 53437 1577 53483
rect 1623 53437 1701 53483
rect 1747 53437 1825 53483
rect 1871 53437 1949 53483
rect 1995 53437 2073 53483
rect 2119 53437 2197 53483
rect 2243 53437 2321 53483
rect 2367 53437 2445 53483
rect 2491 53437 2569 53483
rect 2615 53437 2693 53483
rect 2739 53437 2817 53483
rect 2863 53437 2941 53483
rect 2987 53437 3065 53483
rect 3111 53437 3189 53483
rect 3235 53437 3313 53483
rect 3359 53437 3437 53483
rect 3483 53437 3561 53483
rect 3607 53437 3685 53483
rect 3731 53437 3809 53483
rect 3855 53437 3933 53483
rect 3979 53437 4057 53483
rect 4103 53437 4181 53483
rect 4227 53437 4305 53483
rect 4351 53437 4429 53483
rect 4475 53437 4553 53483
rect 4599 53437 4677 53483
rect 4723 53437 4801 53483
rect 4847 53437 4925 53483
rect 4971 53437 5049 53483
rect 5095 53437 5173 53483
rect 5219 53437 5297 53483
rect 5343 53437 5421 53483
rect 5467 53437 5545 53483
rect 5591 53437 5669 53483
rect 5715 53437 5793 53483
rect 5839 53437 5917 53483
rect 5963 53437 6041 53483
rect 6087 53437 6165 53483
rect 6211 53437 6289 53483
rect 6335 53437 6413 53483
rect 6459 53437 6537 53483
rect 6583 53437 6661 53483
rect 6707 53437 6785 53483
rect 6831 53437 6909 53483
rect 6955 53437 7033 53483
rect 7079 53437 7157 53483
rect 7203 53437 7281 53483
rect 7327 53437 7405 53483
rect 7451 53437 7529 53483
rect 7575 53437 7653 53483
rect 7699 53437 7777 53483
rect 7823 53437 7901 53483
rect 7947 53437 8025 53483
rect 8071 53437 8149 53483
rect 8195 53437 8273 53483
rect 8319 53437 8397 53483
rect 8443 53437 8521 53483
rect 8567 53437 8645 53483
rect 8691 53437 8769 53483
rect 8815 53437 8893 53483
rect 8939 53437 9017 53483
rect 9063 53437 9141 53483
rect 9187 53437 9265 53483
rect 9311 53437 9389 53483
rect 9435 53437 9513 53483
rect 9559 53437 9637 53483
rect 9683 53437 9761 53483
rect 9807 53437 9885 53483
rect 9931 53437 10009 53483
rect 10055 53437 10133 53483
rect 10179 53437 10257 53483
rect 10303 53437 10381 53483
rect 10427 53437 10505 53483
rect 10551 53437 10629 53483
rect 10675 53437 10753 53483
rect 10799 53437 10877 53483
rect 10923 53437 11001 53483
rect 11047 53437 11125 53483
rect 11171 53437 11249 53483
rect 11295 53437 11373 53483
rect 11419 53437 11497 53483
rect 11543 53437 11621 53483
rect 11667 53437 11745 53483
rect 11791 53437 11869 53483
rect 11915 53437 11993 53483
rect 12039 53437 12117 53483
rect 12163 53437 12241 53483
rect 12287 53437 12365 53483
rect 12411 53437 12489 53483
rect 12535 53437 12613 53483
rect 12659 53437 12737 53483
rect 12783 53437 12861 53483
rect 12907 53437 12985 53483
rect 13031 53437 13109 53483
rect 13155 53437 13233 53483
rect 13279 53437 13357 53483
rect 13403 53437 13481 53483
rect 13527 53437 13605 53483
rect 13651 53437 13729 53483
rect 13775 53437 13853 53483
rect 13899 53437 13977 53483
rect 14023 53437 14101 53483
rect 14147 53437 14225 53483
rect 14271 53437 14349 53483
rect 14395 53437 14473 53483
rect 14519 53437 14597 53483
rect 14643 53437 14721 53483
rect 14767 53437 14845 53483
rect 14891 53437 14969 53483
rect 15015 53437 15093 53483
rect 15139 53437 15217 53483
rect 15263 53437 15341 53483
rect 15387 53437 15465 53483
rect 15511 53437 15589 53483
rect 15635 53437 15713 53483
rect 15759 53437 15837 53483
rect 15883 53437 15961 53483
rect 16007 53437 16085 53483
rect 16131 53437 16209 53483
rect 16255 53437 16333 53483
rect 16379 53437 16457 53483
rect 16503 53437 16581 53483
rect 16627 53437 16705 53483
rect 16751 53437 16829 53483
rect 16875 53437 16953 53483
rect 16999 53437 17077 53483
rect 17123 53437 17201 53483
rect 17247 53437 17325 53483
rect 17371 53437 17449 53483
rect 17495 53437 17573 53483
rect 17619 53437 17697 53483
rect 17743 53437 17821 53483
rect 17867 53437 17945 53483
rect 17991 53437 18069 53483
rect 18115 53437 18193 53483
rect 18239 53437 18317 53483
rect 18363 53437 18441 53483
rect 18487 53437 18565 53483
rect 18611 53437 18689 53483
rect 18735 53437 18813 53483
rect 18859 53437 18937 53483
rect 18983 53437 19061 53483
rect 19107 53437 19185 53483
rect 19231 53437 19309 53483
rect 19355 53437 19433 53483
rect 19479 53437 19557 53483
rect 19603 53437 19681 53483
rect 19727 53437 19805 53483
rect 19851 53437 19929 53483
rect 19975 53437 20053 53483
rect 20099 53437 20177 53483
rect 20223 53437 20301 53483
rect 20347 53437 20425 53483
rect 20471 53437 20549 53483
rect 20595 53437 20673 53483
rect 20719 53437 20797 53483
rect 20843 53437 20921 53483
rect 20967 53437 21045 53483
rect 21091 53437 21169 53483
rect 21215 53437 21293 53483
rect 21339 53437 21417 53483
rect 21463 53437 21541 53483
rect 21587 53437 21665 53483
rect 21711 53437 21789 53483
rect 21835 53437 21913 53483
rect 21959 53437 22037 53483
rect 22083 53437 22161 53483
rect 22207 53437 22285 53483
rect 22331 53437 22409 53483
rect 22455 53437 22533 53483
rect 22579 53437 22657 53483
rect 22703 53437 22781 53483
rect 22827 53437 22905 53483
rect 22951 53437 23029 53483
rect 23075 53437 23153 53483
rect 23199 53437 23277 53483
rect 23323 53437 23401 53483
rect 23447 53437 23525 53483
rect 23571 53437 23649 53483
rect 23695 53437 23773 53483
rect 23819 53437 23897 53483
rect 23943 53437 24021 53483
rect 24067 53437 24145 53483
rect 24191 53437 24269 53483
rect 24315 53437 24393 53483
rect 24439 53437 24517 53483
rect 24563 53437 24641 53483
rect 24687 53437 24765 53483
rect 24811 53437 24889 53483
rect 24935 53437 25013 53483
rect 25059 53437 25137 53483
rect 25183 53437 25261 53483
rect 25307 53437 25385 53483
rect 25431 53437 25509 53483
rect 25555 53437 25633 53483
rect 25679 53437 25757 53483
rect 25803 53437 25881 53483
rect 25927 53437 26005 53483
rect 26051 53437 26129 53483
rect 26175 53437 26253 53483
rect 26299 53437 26377 53483
rect 26423 53437 26501 53483
rect 26547 53437 26625 53483
rect 26671 53437 26749 53483
rect 26795 53437 26873 53483
rect 26919 53437 26997 53483
rect 27043 53437 27121 53483
rect 27167 53437 27245 53483
rect 27291 53437 27369 53483
rect 27415 53437 27493 53483
rect 27539 53437 27617 53483
rect 27663 53437 27741 53483
rect 27787 53437 27865 53483
rect 27911 53437 27989 53483
rect 28035 53437 28113 53483
rect 28159 53437 28237 53483
rect 28283 53437 28361 53483
rect 28407 53437 28485 53483
rect 28531 53437 28609 53483
rect 28655 53437 28733 53483
rect 28779 53437 28857 53483
rect 28903 53437 28981 53483
rect 29027 53437 29105 53483
rect 29151 53437 29229 53483
rect 29275 53437 29353 53483
rect 29399 53437 29477 53483
rect 29523 53437 29601 53483
rect 29647 53437 29725 53483
rect 29771 53437 29849 53483
rect 29895 53437 29973 53483
rect 30019 53437 30097 53483
rect 30143 53437 30221 53483
rect 30267 53437 30345 53483
rect 30391 53437 30469 53483
rect 30515 53437 30593 53483
rect 30639 53437 30717 53483
rect 30763 53437 30841 53483
rect 30887 53437 30965 53483
rect 31011 53437 31089 53483
rect 31135 53437 31213 53483
rect 31259 53437 31337 53483
rect 31383 53437 31461 53483
rect 31507 53437 31585 53483
rect 31631 53437 31709 53483
rect 31755 53437 31833 53483
rect 31879 53437 31957 53483
rect 32003 53437 32081 53483
rect 32127 53437 32205 53483
rect 32251 53437 32329 53483
rect 32375 53437 32453 53483
rect 32499 53437 32577 53483
rect 32623 53437 32701 53483
rect 32747 53437 32825 53483
rect 32871 53437 32949 53483
rect 32995 53437 33073 53483
rect 33119 53437 33197 53483
rect 33243 53437 33321 53483
rect 33367 53437 33445 53483
rect 33491 53437 33569 53483
rect 33615 53437 33693 53483
rect 33739 53437 33817 53483
rect 33863 53437 33941 53483
rect 33987 53437 34065 53483
rect 34111 53437 34189 53483
rect 34235 53437 34313 53483
rect 34359 53437 34437 53483
rect 34483 53437 34561 53483
rect 34607 53437 34685 53483
rect 34731 53437 34809 53483
rect 34855 53437 34933 53483
rect 34979 53437 35057 53483
rect 35103 53437 35181 53483
rect 35227 53437 35305 53483
rect 35351 53437 35429 53483
rect 35475 53437 35553 53483
rect 35599 53437 35677 53483
rect 35723 53437 35801 53483
rect 35847 53437 35925 53483
rect 35971 53437 36049 53483
rect 36095 53437 36173 53483
rect 36219 53437 36297 53483
rect 36343 53437 36421 53483
rect 36467 53437 36545 53483
rect 36591 53437 36669 53483
rect 36715 53437 36793 53483
rect 36839 53437 36917 53483
rect 36963 53437 37041 53483
rect 37087 53437 37165 53483
rect 37211 53437 37289 53483
rect 37335 53437 37413 53483
rect 37459 53437 37537 53483
rect 37583 53437 37661 53483
rect 37707 53437 37785 53483
rect 37831 53437 37909 53483
rect 37955 53437 38033 53483
rect 38079 53437 38157 53483
rect 38203 53437 38281 53483
rect 38327 53437 38405 53483
rect 38451 53437 38529 53483
rect 38575 53437 38653 53483
rect 38699 53437 38777 53483
rect 38823 53437 38901 53483
rect 38947 53437 39025 53483
rect 39071 53437 39149 53483
rect 39195 53437 39273 53483
rect 39319 53437 39397 53483
rect 39443 53437 39521 53483
rect 39567 53437 39645 53483
rect 39691 53437 39769 53483
rect 39815 53437 39893 53483
rect 39939 53437 40017 53483
rect 40063 53437 40141 53483
rect 40187 53437 40265 53483
rect 40311 53437 40389 53483
rect 40435 53437 40513 53483
rect 40559 53437 40637 53483
rect 40683 53437 40761 53483
rect 40807 53437 40885 53483
rect 40931 53437 41009 53483
rect 41055 53437 41133 53483
rect 41179 53437 41257 53483
rect 41303 53437 41381 53483
rect 41427 53437 41505 53483
rect 41551 53437 41629 53483
rect 41675 53437 41753 53483
rect 41799 53437 41877 53483
rect 41923 53437 42001 53483
rect 42047 53437 42125 53483
rect 42171 53437 42249 53483
rect 42295 53437 42373 53483
rect 42419 53437 42497 53483
rect 42543 53437 42621 53483
rect 42667 53437 42745 53483
rect 42791 53437 42869 53483
rect 42915 53437 42993 53483
rect 43039 53437 43117 53483
rect 43163 53437 43241 53483
rect 43287 53437 43365 53483
rect 43411 53437 43489 53483
rect 43535 53437 43613 53483
rect 43659 53437 43737 53483
rect 43783 53437 43861 53483
rect 43907 53437 43985 53483
rect 44031 53437 44109 53483
rect 44155 53437 44233 53483
rect 44279 53437 44357 53483
rect 44403 53437 44481 53483
rect 44527 53437 44605 53483
rect 44651 53437 44729 53483
rect 44775 53437 44853 53483
rect 44899 53437 44977 53483
rect 45023 53437 45101 53483
rect 45147 53437 45225 53483
rect 45271 53437 45349 53483
rect 45395 53437 45473 53483
rect 45519 53437 45597 53483
rect 45643 53437 45721 53483
rect 45767 53437 45845 53483
rect 45891 53437 45969 53483
rect 46015 53437 46093 53483
rect 46139 53437 46217 53483
rect 46263 53437 46341 53483
rect 46387 53437 46465 53483
rect 46511 53437 46589 53483
rect 46635 53437 46713 53483
rect 46759 53437 46837 53483
rect 46883 53437 46961 53483
rect 47007 53437 47085 53483
rect 47131 53437 47209 53483
rect 47255 53437 47333 53483
rect 47379 53437 47457 53483
rect 47503 53437 47581 53483
rect 47627 53437 47705 53483
rect 47751 53437 47829 53483
rect 47875 53437 47953 53483
rect 47999 53437 48077 53483
rect 48123 53437 48201 53483
rect 48247 53437 48325 53483
rect 48371 53437 48449 53483
rect 48495 53437 48573 53483
rect 48619 53437 48697 53483
rect 48743 53437 48821 53483
rect 48867 53437 48945 53483
rect 48991 53437 49069 53483
rect 49115 53437 49193 53483
rect 49239 53437 49317 53483
rect 49363 53437 49441 53483
rect 49487 53437 49565 53483
rect 49611 53437 49689 53483
rect 49735 53437 49813 53483
rect 49859 53437 49937 53483
rect 49983 53437 50061 53483
rect 50107 53437 50185 53483
rect 50231 53437 50309 53483
rect 50355 53437 50433 53483
rect 50479 53437 50557 53483
rect 50603 53437 50681 53483
rect 50727 53437 50805 53483
rect 50851 53437 50929 53483
rect 50975 53437 51053 53483
rect 51099 53437 51177 53483
rect 51223 53437 51301 53483
rect 51347 53437 51425 53483
rect 51471 53437 51549 53483
rect 51595 53437 51673 53483
rect 51719 53437 51797 53483
rect 51843 53437 51921 53483
rect 51967 53437 52045 53483
rect 52091 53437 52169 53483
rect 52215 53437 52293 53483
rect 52339 53437 52417 53483
rect 52463 53437 52541 53483
rect 52587 53437 52665 53483
rect 52711 53437 52789 53483
rect 52835 53437 52913 53483
rect 52959 53437 53037 53483
rect 53083 53437 53161 53483
rect 53207 53437 53285 53483
rect 53331 53437 53409 53483
rect 53455 53437 53533 53483
rect 53579 53437 53657 53483
rect 53703 53437 53781 53483
rect 53827 53437 53905 53483
rect 53951 53437 54029 53483
rect 54075 53437 54153 53483
rect 54199 53437 54277 53483
rect 54323 53437 54401 53483
rect 54447 53437 54525 53483
rect 54571 53437 54649 53483
rect 54695 53437 54773 53483
rect 54819 53437 54897 53483
rect 54943 53437 55021 53483
rect 55067 53437 55145 53483
rect 55191 53437 55269 53483
rect 55315 53437 55393 53483
rect 55439 53437 55517 53483
rect 55563 53437 55641 53483
rect 55687 53437 55765 53483
rect 55811 53437 55889 53483
rect 55935 53437 56013 53483
rect 56059 53437 56137 53483
rect 56183 53437 56261 53483
rect 56307 53437 56385 53483
rect 56431 53437 56509 53483
rect 56555 53437 56633 53483
rect 56679 53437 56757 53483
rect 56803 53437 56881 53483
rect 56927 53437 57005 53483
rect 57051 53437 57129 53483
rect 57175 53437 57253 53483
rect 57299 53437 57377 53483
rect 57423 53437 57501 53483
rect 57547 53437 57625 53483
rect 57671 53437 57749 53483
rect 57795 53437 57873 53483
rect 57919 53437 57997 53483
rect 58043 53437 58121 53483
rect 58167 53437 58245 53483
rect 58291 53437 58369 53483
rect 58415 53437 58493 53483
rect 58539 53437 58617 53483
rect 58663 53437 58741 53483
rect 58787 53437 58865 53483
rect 58911 53437 58989 53483
rect 59035 53437 59113 53483
rect 59159 53437 59237 53483
rect 59283 53437 59361 53483
rect 59407 53437 59485 53483
rect 59531 53437 59609 53483
rect 59655 53437 59733 53483
rect 59779 53437 59857 53483
rect 59903 53437 59981 53483
rect 60027 53437 60105 53483
rect 60151 53437 60229 53483
rect 60275 53437 60353 53483
rect 60399 53437 60477 53483
rect 60523 53437 60601 53483
rect 60647 53437 60725 53483
rect 60771 53437 60849 53483
rect 60895 53437 60973 53483
rect 61019 53437 61097 53483
rect 61143 53437 61221 53483
rect 61267 53437 61345 53483
rect 61391 53437 61469 53483
rect 61515 53437 61593 53483
rect 61639 53437 61717 53483
rect 61763 53437 61841 53483
rect 61887 53437 61965 53483
rect 62011 53437 62089 53483
rect 62135 53437 62213 53483
rect 62259 53437 62337 53483
rect 62383 53437 62461 53483
rect 62507 53437 62585 53483
rect 62631 53437 62709 53483
rect 62755 53437 62833 53483
rect 62879 53437 62957 53483
rect 63003 53437 63081 53483
rect 63127 53437 63205 53483
rect 63251 53437 63329 53483
rect 63375 53437 63453 53483
rect 63499 53437 63577 53483
rect 63623 53437 63701 53483
rect 63747 53437 63825 53483
rect 63871 53437 63949 53483
rect 63995 53437 64073 53483
rect 64119 53437 64197 53483
rect 64243 53437 64321 53483
rect 64367 53437 64445 53483
rect 64491 53437 64569 53483
rect 64615 53437 64693 53483
rect 64739 53437 64817 53483
rect 64863 53437 64941 53483
rect 64987 53437 65065 53483
rect 65111 53437 65189 53483
rect 65235 53437 65313 53483
rect 65359 53437 65437 53483
rect 65483 53437 65561 53483
rect 65607 53437 65685 53483
rect 65731 53437 65809 53483
rect 65855 53437 65933 53483
rect 65979 53437 66057 53483
rect 66103 53437 66181 53483
rect 66227 53437 66305 53483
rect 66351 53437 66429 53483
rect 66475 53437 66553 53483
rect 66599 53437 66677 53483
rect 66723 53437 66801 53483
rect 66847 53437 66925 53483
rect 66971 53437 67049 53483
rect 67095 53437 67173 53483
rect 67219 53437 67297 53483
rect 67343 53437 67421 53483
rect 67467 53437 67545 53483
rect 67591 53437 67669 53483
rect 67715 53437 67793 53483
rect 67839 53437 67917 53483
rect 67963 53437 68041 53483
rect 68087 53437 68165 53483
rect 68211 53437 68289 53483
rect 68335 53437 68413 53483
rect 68459 53437 68537 53483
rect 68583 53437 68661 53483
rect 68707 53437 68785 53483
rect 68831 53437 68909 53483
rect 68955 53437 69033 53483
rect 69079 53437 69157 53483
rect 69203 53437 69281 53483
rect 69327 53437 69405 53483
rect 69451 53437 69529 53483
rect 69575 53437 69653 53483
rect 69699 53437 69777 53483
rect 69823 53437 69901 53483
rect 69947 53437 70025 53483
rect 70071 53437 70149 53483
rect 70195 53437 70273 53483
rect 70319 53437 70397 53483
rect 70443 53437 70521 53483
rect 70567 53437 70645 53483
rect 70691 53437 70769 53483
rect 70815 53437 70893 53483
rect 70939 53437 71017 53483
rect 71063 53437 71141 53483
rect 71187 53437 71265 53483
rect 71311 53437 71389 53483
rect 71435 53437 71513 53483
rect 71559 53437 71637 53483
rect 71683 53437 71761 53483
rect 71807 53437 71885 53483
rect 71931 53437 72009 53483
rect 72055 53437 72133 53483
rect 72179 53437 72257 53483
rect 72303 53437 72381 53483
rect 72427 53437 72505 53483
rect 72551 53437 72629 53483
rect 72675 53437 72753 53483
rect 72799 53437 72877 53483
rect 72923 53437 73001 53483
rect 73047 53437 73125 53483
rect 73171 53437 73249 53483
rect 73295 53437 73373 53483
rect 73419 53437 73497 53483
rect 73543 53437 73621 53483
rect 73667 53437 73745 53483
rect 73791 53437 73869 53483
rect 73915 53437 73993 53483
rect 74039 53437 74117 53483
rect 74163 53437 74241 53483
rect 74287 53437 74365 53483
rect 74411 53437 74489 53483
rect 74535 53437 74613 53483
rect 74659 53437 74737 53483
rect 74783 53437 74861 53483
rect 74907 53437 74985 53483
rect 75031 53437 75109 53483
rect 75155 53437 75233 53483
rect 75279 53437 75357 53483
rect 75403 53437 75481 53483
rect 75527 53437 75605 53483
rect 75651 53437 75729 53483
rect 75775 53437 75853 53483
rect 75899 53437 75977 53483
rect 76023 53437 76101 53483
rect 76147 53437 76225 53483
rect 76271 53437 76349 53483
rect 76395 53437 76473 53483
rect 76519 53437 76597 53483
rect 76643 53437 76721 53483
rect 76767 53437 76845 53483
rect 76891 53437 76969 53483
rect 77015 53437 77093 53483
rect 77139 53437 77217 53483
rect 77263 53437 77341 53483
rect 77387 53437 77465 53483
rect 77511 53437 77589 53483
rect 77635 53437 77713 53483
rect 77759 53437 77837 53483
rect 77883 53437 77961 53483
rect 78007 53437 78085 53483
rect 78131 53437 78209 53483
rect 78255 53437 78333 53483
rect 78379 53437 78457 53483
rect 78503 53437 78581 53483
rect 78627 53437 78705 53483
rect 78751 53437 78829 53483
rect 78875 53437 78953 53483
rect 78999 53437 79077 53483
rect 79123 53437 79201 53483
rect 79247 53437 79325 53483
rect 79371 53437 79449 53483
rect 79495 53437 79573 53483
rect 79619 53437 79697 53483
rect 79743 53437 79821 53483
rect 79867 53437 79945 53483
rect 79991 53437 80069 53483
rect 80115 53437 80193 53483
rect 80239 53437 80317 53483
rect 80363 53437 80441 53483
rect 80487 53437 80565 53483
rect 80611 53437 80689 53483
rect 80735 53437 80813 53483
rect 80859 53437 80937 53483
rect 80983 53437 81061 53483
rect 81107 53437 81185 53483
rect 81231 53437 81309 53483
rect 81355 53437 81433 53483
rect 81479 53437 81557 53483
rect 81603 53437 81681 53483
rect 81727 53437 81805 53483
rect 81851 53437 81929 53483
rect 81975 53437 82053 53483
rect 82099 53437 82177 53483
rect 82223 53437 82301 53483
rect 82347 53437 82425 53483
rect 82471 53437 82549 53483
rect 82595 53437 82673 53483
rect 82719 53437 82797 53483
rect 82843 53437 82921 53483
rect 82967 53437 83045 53483
rect 83091 53437 83169 53483
rect 83215 53437 83293 53483
rect 83339 53437 83417 53483
rect 83463 53437 83541 53483
rect 83587 53437 83665 53483
rect 83711 53437 83789 53483
rect 83835 53437 83913 53483
rect 83959 53437 84037 53483
rect 84083 53437 84161 53483
rect 84207 53437 84285 53483
rect 84331 53437 84409 53483
rect 84455 53437 84533 53483
rect 84579 53437 84657 53483
rect 84703 53437 84781 53483
rect 84827 53437 84905 53483
rect 84951 53437 85029 53483
rect 85075 53437 85153 53483
rect 85199 53437 85277 53483
rect 85323 53437 85401 53483
rect 85447 53437 85525 53483
rect 85571 53437 85649 53483
rect 85695 53437 85706 53483
rect 0 53359 85706 53437
rect 0 53313 89 53359
rect 135 53313 213 53359
rect 259 53313 337 53359
rect 383 53313 461 53359
rect 507 53313 585 53359
rect 631 53313 709 53359
rect 755 53313 833 53359
rect 879 53313 957 53359
rect 1003 53313 1081 53359
rect 1127 53313 1205 53359
rect 1251 53313 1329 53359
rect 1375 53313 1453 53359
rect 1499 53313 1577 53359
rect 1623 53313 1701 53359
rect 1747 53313 1825 53359
rect 1871 53313 1949 53359
rect 1995 53313 2073 53359
rect 2119 53313 2197 53359
rect 2243 53313 2321 53359
rect 2367 53313 2445 53359
rect 2491 53313 2569 53359
rect 2615 53313 2693 53359
rect 2739 53313 2817 53359
rect 2863 53313 2941 53359
rect 2987 53313 3065 53359
rect 3111 53313 3189 53359
rect 3235 53313 3313 53359
rect 3359 53313 3437 53359
rect 3483 53313 3561 53359
rect 3607 53313 3685 53359
rect 3731 53313 3809 53359
rect 3855 53313 3933 53359
rect 3979 53313 4057 53359
rect 4103 53313 4181 53359
rect 4227 53313 4305 53359
rect 4351 53313 4429 53359
rect 4475 53313 4553 53359
rect 4599 53313 4677 53359
rect 4723 53313 4801 53359
rect 4847 53313 4925 53359
rect 4971 53313 5049 53359
rect 5095 53313 5173 53359
rect 5219 53313 5297 53359
rect 5343 53313 5421 53359
rect 5467 53313 5545 53359
rect 5591 53313 5669 53359
rect 5715 53313 5793 53359
rect 5839 53313 5917 53359
rect 5963 53313 6041 53359
rect 6087 53313 6165 53359
rect 6211 53313 6289 53359
rect 6335 53313 6413 53359
rect 6459 53313 6537 53359
rect 6583 53313 6661 53359
rect 6707 53313 6785 53359
rect 6831 53313 6909 53359
rect 6955 53313 7033 53359
rect 7079 53313 7157 53359
rect 7203 53313 7281 53359
rect 7327 53313 7405 53359
rect 7451 53313 7529 53359
rect 7575 53313 7653 53359
rect 7699 53313 7777 53359
rect 7823 53313 7901 53359
rect 7947 53313 8025 53359
rect 8071 53313 8149 53359
rect 8195 53313 8273 53359
rect 8319 53313 8397 53359
rect 8443 53313 8521 53359
rect 8567 53313 8645 53359
rect 8691 53313 8769 53359
rect 8815 53313 8893 53359
rect 8939 53313 9017 53359
rect 9063 53313 9141 53359
rect 9187 53313 9265 53359
rect 9311 53313 9389 53359
rect 9435 53313 9513 53359
rect 9559 53313 9637 53359
rect 9683 53313 9761 53359
rect 9807 53313 9885 53359
rect 9931 53313 10009 53359
rect 10055 53313 10133 53359
rect 10179 53313 10257 53359
rect 10303 53313 10381 53359
rect 10427 53313 10505 53359
rect 10551 53313 10629 53359
rect 10675 53313 10753 53359
rect 10799 53313 10877 53359
rect 10923 53313 11001 53359
rect 11047 53313 11125 53359
rect 11171 53313 11249 53359
rect 11295 53313 11373 53359
rect 11419 53313 11497 53359
rect 11543 53313 11621 53359
rect 11667 53313 11745 53359
rect 11791 53313 11869 53359
rect 11915 53313 11993 53359
rect 12039 53313 12117 53359
rect 12163 53313 12241 53359
rect 12287 53313 12365 53359
rect 12411 53313 12489 53359
rect 12535 53313 12613 53359
rect 12659 53313 12737 53359
rect 12783 53313 12861 53359
rect 12907 53313 12985 53359
rect 13031 53313 13109 53359
rect 13155 53313 13233 53359
rect 13279 53313 13357 53359
rect 13403 53313 13481 53359
rect 13527 53313 13605 53359
rect 13651 53313 13729 53359
rect 13775 53313 13853 53359
rect 13899 53313 13977 53359
rect 14023 53313 14101 53359
rect 14147 53313 14225 53359
rect 14271 53313 14349 53359
rect 14395 53313 14473 53359
rect 14519 53313 14597 53359
rect 14643 53313 14721 53359
rect 14767 53313 14845 53359
rect 14891 53313 14969 53359
rect 15015 53313 15093 53359
rect 15139 53313 15217 53359
rect 15263 53313 15341 53359
rect 15387 53313 15465 53359
rect 15511 53313 15589 53359
rect 15635 53313 15713 53359
rect 15759 53313 15837 53359
rect 15883 53313 15961 53359
rect 16007 53313 16085 53359
rect 16131 53313 16209 53359
rect 16255 53313 16333 53359
rect 16379 53313 16457 53359
rect 16503 53313 16581 53359
rect 16627 53313 16705 53359
rect 16751 53313 16829 53359
rect 16875 53313 16953 53359
rect 16999 53313 17077 53359
rect 17123 53313 17201 53359
rect 17247 53313 17325 53359
rect 17371 53313 17449 53359
rect 17495 53313 17573 53359
rect 17619 53313 17697 53359
rect 17743 53313 17821 53359
rect 17867 53313 17945 53359
rect 17991 53313 18069 53359
rect 18115 53313 18193 53359
rect 18239 53313 18317 53359
rect 18363 53313 18441 53359
rect 18487 53313 18565 53359
rect 18611 53313 18689 53359
rect 18735 53313 18813 53359
rect 18859 53313 18937 53359
rect 18983 53313 19061 53359
rect 19107 53313 19185 53359
rect 19231 53313 19309 53359
rect 19355 53313 19433 53359
rect 19479 53313 19557 53359
rect 19603 53313 19681 53359
rect 19727 53313 19805 53359
rect 19851 53313 19929 53359
rect 19975 53313 20053 53359
rect 20099 53313 20177 53359
rect 20223 53313 20301 53359
rect 20347 53313 20425 53359
rect 20471 53313 20549 53359
rect 20595 53313 20673 53359
rect 20719 53313 20797 53359
rect 20843 53313 20921 53359
rect 20967 53313 21045 53359
rect 21091 53313 21169 53359
rect 21215 53313 21293 53359
rect 21339 53313 21417 53359
rect 21463 53313 21541 53359
rect 21587 53313 21665 53359
rect 21711 53313 21789 53359
rect 21835 53313 21913 53359
rect 21959 53313 22037 53359
rect 22083 53313 22161 53359
rect 22207 53313 22285 53359
rect 22331 53313 22409 53359
rect 22455 53313 22533 53359
rect 22579 53313 22657 53359
rect 22703 53313 22781 53359
rect 22827 53313 22905 53359
rect 22951 53313 23029 53359
rect 23075 53313 23153 53359
rect 23199 53313 23277 53359
rect 23323 53313 23401 53359
rect 23447 53313 23525 53359
rect 23571 53313 23649 53359
rect 23695 53313 23773 53359
rect 23819 53313 23897 53359
rect 23943 53313 24021 53359
rect 24067 53313 24145 53359
rect 24191 53313 24269 53359
rect 24315 53313 24393 53359
rect 24439 53313 24517 53359
rect 24563 53313 24641 53359
rect 24687 53313 24765 53359
rect 24811 53313 24889 53359
rect 24935 53313 25013 53359
rect 25059 53313 25137 53359
rect 25183 53313 25261 53359
rect 25307 53313 25385 53359
rect 25431 53313 25509 53359
rect 25555 53313 25633 53359
rect 25679 53313 25757 53359
rect 25803 53313 25881 53359
rect 25927 53313 26005 53359
rect 26051 53313 26129 53359
rect 26175 53313 26253 53359
rect 26299 53313 26377 53359
rect 26423 53313 26501 53359
rect 26547 53313 26625 53359
rect 26671 53313 26749 53359
rect 26795 53313 26873 53359
rect 26919 53313 26997 53359
rect 27043 53313 27121 53359
rect 27167 53313 27245 53359
rect 27291 53313 27369 53359
rect 27415 53313 27493 53359
rect 27539 53313 27617 53359
rect 27663 53313 27741 53359
rect 27787 53313 27865 53359
rect 27911 53313 27989 53359
rect 28035 53313 28113 53359
rect 28159 53313 28237 53359
rect 28283 53313 28361 53359
rect 28407 53313 28485 53359
rect 28531 53313 28609 53359
rect 28655 53313 28733 53359
rect 28779 53313 28857 53359
rect 28903 53313 28981 53359
rect 29027 53313 29105 53359
rect 29151 53313 29229 53359
rect 29275 53313 29353 53359
rect 29399 53313 29477 53359
rect 29523 53313 29601 53359
rect 29647 53313 29725 53359
rect 29771 53313 29849 53359
rect 29895 53313 29973 53359
rect 30019 53313 30097 53359
rect 30143 53313 30221 53359
rect 30267 53313 30345 53359
rect 30391 53313 30469 53359
rect 30515 53313 30593 53359
rect 30639 53313 30717 53359
rect 30763 53313 30841 53359
rect 30887 53313 30965 53359
rect 31011 53313 31089 53359
rect 31135 53313 31213 53359
rect 31259 53313 31337 53359
rect 31383 53313 31461 53359
rect 31507 53313 31585 53359
rect 31631 53313 31709 53359
rect 31755 53313 31833 53359
rect 31879 53313 31957 53359
rect 32003 53313 32081 53359
rect 32127 53313 32205 53359
rect 32251 53313 32329 53359
rect 32375 53313 32453 53359
rect 32499 53313 32577 53359
rect 32623 53313 32701 53359
rect 32747 53313 32825 53359
rect 32871 53313 32949 53359
rect 32995 53313 33073 53359
rect 33119 53313 33197 53359
rect 33243 53313 33321 53359
rect 33367 53313 33445 53359
rect 33491 53313 33569 53359
rect 33615 53313 33693 53359
rect 33739 53313 33817 53359
rect 33863 53313 33941 53359
rect 33987 53313 34065 53359
rect 34111 53313 34189 53359
rect 34235 53313 34313 53359
rect 34359 53313 34437 53359
rect 34483 53313 34561 53359
rect 34607 53313 34685 53359
rect 34731 53313 34809 53359
rect 34855 53313 34933 53359
rect 34979 53313 35057 53359
rect 35103 53313 35181 53359
rect 35227 53313 35305 53359
rect 35351 53313 35429 53359
rect 35475 53313 35553 53359
rect 35599 53313 35677 53359
rect 35723 53313 35801 53359
rect 35847 53313 35925 53359
rect 35971 53313 36049 53359
rect 36095 53313 36173 53359
rect 36219 53313 36297 53359
rect 36343 53313 36421 53359
rect 36467 53313 36545 53359
rect 36591 53313 36669 53359
rect 36715 53313 36793 53359
rect 36839 53313 36917 53359
rect 36963 53313 37041 53359
rect 37087 53313 37165 53359
rect 37211 53313 37289 53359
rect 37335 53313 37413 53359
rect 37459 53313 37537 53359
rect 37583 53313 37661 53359
rect 37707 53313 37785 53359
rect 37831 53313 37909 53359
rect 37955 53313 38033 53359
rect 38079 53313 38157 53359
rect 38203 53313 38281 53359
rect 38327 53313 38405 53359
rect 38451 53313 38529 53359
rect 38575 53313 38653 53359
rect 38699 53313 38777 53359
rect 38823 53313 38901 53359
rect 38947 53313 39025 53359
rect 39071 53313 39149 53359
rect 39195 53313 39273 53359
rect 39319 53313 39397 53359
rect 39443 53313 39521 53359
rect 39567 53313 39645 53359
rect 39691 53313 39769 53359
rect 39815 53313 39893 53359
rect 39939 53313 40017 53359
rect 40063 53313 40141 53359
rect 40187 53313 40265 53359
rect 40311 53313 40389 53359
rect 40435 53313 40513 53359
rect 40559 53313 40637 53359
rect 40683 53313 40761 53359
rect 40807 53313 40885 53359
rect 40931 53313 41009 53359
rect 41055 53313 41133 53359
rect 41179 53313 41257 53359
rect 41303 53313 41381 53359
rect 41427 53313 41505 53359
rect 41551 53313 41629 53359
rect 41675 53313 41753 53359
rect 41799 53313 41877 53359
rect 41923 53313 42001 53359
rect 42047 53313 42125 53359
rect 42171 53313 42249 53359
rect 42295 53313 42373 53359
rect 42419 53313 42497 53359
rect 42543 53313 42621 53359
rect 42667 53313 42745 53359
rect 42791 53313 42869 53359
rect 42915 53313 42993 53359
rect 43039 53313 43117 53359
rect 43163 53313 43241 53359
rect 43287 53313 43365 53359
rect 43411 53313 43489 53359
rect 43535 53313 43613 53359
rect 43659 53313 43737 53359
rect 43783 53313 43861 53359
rect 43907 53313 43985 53359
rect 44031 53313 44109 53359
rect 44155 53313 44233 53359
rect 44279 53313 44357 53359
rect 44403 53313 44481 53359
rect 44527 53313 44605 53359
rect 44651 53313 44729 53359
rect 44775 53313 44853 53359
rect 44899 53313 44977 53359
rect 45023 53313 45101 53359
rect 45147 53313 45225 53359
rect 45271 53313 45349 53359
rect 45395 53313 45473 53359
rect 45519 53313 45597 53359
rect 45643 53313 45721 53359
rect 45767 53313 45845 53359
rect 45891 53313 45969 53359
rect 46015 53313 46093 53359
rect 46139 53313 46217 53359
rect 46263 53313 46341 53359
rect 46387 53313 46465 53359
rect 46511 53313 46589 53359
rect 46635 53313 46713 53359
rect 46759 53313 46837 53359
rect 46883 53313 46961 53359
rect 47007 53313 47085 53359
rect 47131 53313 47209 53359
rect 47255 53313 47333 53359
rect 47379 53313 47457 53359
rect 47503 53313 47581 53359
rect 47627 53313 47705 53359
rect 47751 53313 47829 53359
rect 47875 53313 47953 53359
rect 47999 53313 48077 53359
rect 48123 53313 48201 53359
rect 48247 53313 48325 53359
rect 48371 53313 48449 53359
rect 48495 53313 48573 53359
rect 48619 53313 48697 53359
rect 48743 53313 48821 53359
rect 48867 53313 48945 53359
rect 48991 53313 49069 53359
rect 49115 53313 49193 53359
rect 49239 53313 49317 53359
rect 49363 53313 49441 53359
rect 49487 53313 49565 53359
rect 49611 53313 49689 53359
rect 49735 53313 49813 53359
rect 49859 53313 49937 53359
rect 49983 53313 50061 53359
rect 50107 53313 50185 53359
rect 50231 53313 50309 53359
rect 50355 53313 50433 53359
rect 50479 53313 50557 53359
rect 50603 53313 50681 53359
rect 50727 53313 50805 53359
rect 50851 53313 50929 53359
rect 50975 53313 51053 53359
rect 51099 53313 51177 53359
rect 51223 53313 51301 53359
rect 51347 53313 51425 53359
rect 51471 53313 51549 53359
rect 51595 53313 51673 53359
rect 51719 53313 51797 53359
rect 51843 53313 51921 53359
rect 51967 53313 52045 53359
rect 52091 53313 52169 53359
rect 52215 53313 52293 53359
rect 52339 53313 52417 53359
rect 52463 53313 52541 53359
rect 52587 53313 52665 53359
rect 52711 53313 52789 53359
rect 52835 53313 52913 53359
rect 52959 53313 53037 53359
rect 53083 53313 53161 53359
rect 53207 53313 53285 53359
rect 53331 53313 53409 53359
rect 53455 53313 53533 53359
rect 53579 53313 53657 53359
rect 53703 53313 53781 53359
rect 53827 53313 53905 53359
rect 53951 53313 54029 53359
rect 54075 53313 54153 53359
rect 54199 53313 54277 53359
rect 54323 53313 54401 53359
rect 54447 53313 54525 53359
rect 54571 53313 54649 53359
rect 54695 53313 54773 53359
rect 54819 53313 54897 53359
rect 54943 53313 55021 53359
rect 55067 53313 55145 53359
rect 55191 53313 55269 53359
rect 55315 53313 55393 53359
rect 55439 53313 55517 53359
rect 55563 53313 55641 53359
rect 55687 53313 55765 53359
rect 55811 53313 55889 53359
rect 55935 53313 56013 53359
rect 56059 53313 56137 53359
rect 56183 53313 56261 53359
rect 56307 53313 56385 53359
rect 56431 53313 56509 53359
rect 56555 53313 56633 53359
rect 56679 53313 56757 53359
rect 56803 53313 56881 53359
rect 56927 53313 57005 53359
rect 57051 53313 57129 53359
rect 57175 53313 57253 53359
rect 57299 53313 57377 53359
rect 57423 53313 57501 53359
rect 57547 53313 57625 53359
rect 57671 53313 57749 53359
rect 57795 53313 57873 53359
rect 57919 53313 57997 53359
rect 58043 53313 58121 53359
rect 58167 53313 58245 53359
rect 58291 53313 58369 53359
rect 58415 53313 58493 53359
rect 58539 53313 58617 53359
rect 58663 53313 58741 53359
rect 58787 53313 58865 53359
rect 58911 53313 58989 53359
rect 59035 53313 59113 53359
rect 59159 53313 59237 53359
rect 59283 53313 59361 53359
rect 59407 53313 59485 53359
rect 59531 53313 59609 53359
rect 59655 53313 59733 53359
rect 59779 53313 59857 53359
rect 59903 53313 59981 53359
rect 60027 53313 60105 53359
rect 60151 53313 60229 53359
rect 60275 53313 60353 53359
rect 60399 53313 60477 53359
rect 60523 53313 60601 53359
rect 60647 53313 60725 53359
rect 60771 53313 60849 53359
rect 60895 53313 60973 53359
rect 61019 53313 61097 53359
rect 61143 53313 61221 53359
rect 61267 53313 61345 53359
rect 61391 53313 61469 53359
rect 61515 53313 61593 53359
rect 61639 53313 61717 53359
rect 61763 53313 61841 53359
rect 61887 53313 61965 53359
rect 62011 53313 62089 53359
rect 62135 53313 62213 53359
rect 62259 53313 62337 53359
rect 62383 53313 62461 53359
rect 62507 53313 62585 53359
rect 62631 53313 62709 53359
rect 62755 53313 62833 53359
rect 62879 53313 62957 53359
rect 63003 53313 63081 53359
rect 63127 53313 63205 53359
rect 63251 53313 63329 53359
rect 63375 53313 63453 53359
rect 63499 53313 63577 53359
rect 63623 53313 63701 53359
rect 63747 53313 63825 53359
rect 63871 53313 63949 53359
rect 63995 53313 64073 53359
rect 64119 53313 64197 53359
rect 64243 53313 64321 53359
rect 64367 53313 64445 53359
rect 64491 53313 64569 53359
rect 64615 53313 64693 53359
rect 64739 53313 64817 53359
rect 64863 53313 64941 53359
rect 64987 53313 65065 53359
rect 65111 53313 65189 53359
rect 65235 53313 65313 53359
rect 65359 53313 65437 53359
rect 65483 53313 65561 53359
rect 65607 53313 65685 53359
rect 65731 53313 65809 53359
rect 65855 53313 65933 53359
rect 65979 53313 66057 53359
rect 66103 53313 66181 53359
rect 66227 53313 66305 53359
rect 66351 53313 66429 53359
rect 66475 53313 66553 53359
rect 66599 53313 66677 53359
rect 66723 53313 66801 53359
rect 66847 53313 66925 53359
rect 66971 53313 67049 53359
rect 67095 53313 67173 53359
rect 67219 53313 67297 53359
rect 67343 53313 67421 53359
rect 67467 53313 67545 53359
rect 67591 53313 67669 53359
rect 67715 53313 67793 53359
rect 67839 53313 67917 53359
rect 67963 53313 68041 53359
rect 68087 53313 68165 53359
rect 68211 53313 68289 53359
rect 68335 53313 68413 53359
rect 68459 53313 68537 53359
rect 68583 53313 68661 53359
rect 68707 53313 68785 53359
rect 68831 53313 68909 53359
rect 68955 53313 69033 53359
rect 69079 53313 69157 53359
rect 69203 53313 69281 53359
rect 69327 53313 69405 53359
rect 69451 53313 69529 53359
rect 69575 53313 69653 53359
rect 69699 53313 69777 53359
rect 69823 53313 69901 53359
rect 69947 53313 70025 53359
rect 70071 53313 70149 53359
rect 70195 53313 70273 53359
rect 70319 53313 70397 53359
rect 70443 53313 70521 53359
rect 70567 53313 70645 53359
rect 70691 53313 70769 53359
rect 70815 53313 70893 53359
rect 70939 53313 71017 53359
rect 71063 53313 71141 53359
rect 71187 53313 71265 53359
rect 71311 53313 71389 53359
rect 71435 53313 71513 53359
rect 71559 53313 71637 53359
rect 71683 53313 71761 53359
rect 71807 53313 71885 53359
rect 71931 53313 72009 53359
rect 72055 53313 72133 53359
rect 72179 53313 72257 53359
rect 72303 53313 72381 53359
rect 72427 53313 72505 53359
rect 72551 53313 72629 53359
rect 72675 53313 72753 53359
rect 72799 53313 72877 53359
rect 72923 53313 73001 53359
rect 73047 53313 73125 53359
rect 73171 53313 73249 53359
rect 73295 53313 73373 53359
rect 73419 53313 73497 53359
rect 73543 53313 73621 53359
rect 73667 53313 73745 53359
rect 73791 53313 73869 53359
rect 73915 53313 73993 53359
rect 74039 53313 74117 53359
rect 74163 53313 74241 53359
rect 74287 53313 74365 53359
rect 74411 53313 74489 53359
rect 74535 53313 74613 53359
rect 74659 53313 74737 53359
rect 74783 53313 74861 53359
rect 74907 53313 74985 53359
rect 75031 53313 75109 53359
rect 75155 53313 75233 53359
rect 75279 53313 75357 53359
rect 75403 53313 75481 53359
rect 75527 53313 75605 53359
rect 75651 53313 75729 53359
rect 75775 53313 75853 53359
rect 75899 53313 75977 53359
rect 76023 53313 76101 53359
rect 76147 53313 76225 53359
rect 76271 53313 76349 53359
rect 76395 53313 76473 53359
rect 76519 53313 76597 53359
rect 76643 53313 76721 53359
rect 76767 53313 76845 53359
rect 76891 53313 76969 53359
rect 77015 53313 77093 53359
rect 77139 53313 77217 53359
rect 77263 53313 77341 53359
rect 77387 53313 77465 53359
rect 77511 53313 77589 53359
rect 77635 53313 77713 53359
rect 77759 53313 77837 53359
rect 77883 53313 77961 53359
rect 78007 53313 78085 53359
rect 78131 53313 78209 53359
rect 78255 53313 78333 53359
rect 78379 53313 78457 53359
rect 78503 53313 78581 53359
rect 78627 53313 78705 53359
rect 78751 53313 78829 53359
rect 78875 53313 78953 53359
rect 78999 53313 79077 53359
rect 79123 53313 79201 53359
rect 79247 53313 79325 53359
rect 79371 53313 79449 53359
rect 79495 53313 79573 53359
rect 79619 53313 79697 53359
rect 79743 53313 79821 53359
rect 79867 53313 79945 53359
rect 79991 53313 80069 53359
rect 80115 53313 80193 53359
rect 80239 53313 80317 53359
rect 80363 53313 80441 53359
rect 80487 53313 80565 53359
rect 80611 53313 80689 53359
rect 80735 53313 80813 53359
rect 80859 53313 80937 53359
rect 80983 53313 81061 53359
rect 81107 53313 81185 53359
rect 81231 53313 81309 53359
rect 81355 53313 81433 53359
rect 81479 53313 81557 53359
rect 81603 53313 81681 53359
rect 81727 53313 81805 53359
rect 81851 53313 81929 53359
rect 81975 53313 82053 53359
rect 82099 53313 82177 53359
rect 82223 53313 82301 53359
rect 82347 53313 82425 53359
rect 82471 53313 82549 53359
rect 82595 53313 82673 53359
rect 82719 53313 82797 53359
rect 82843 53313 82921 53359
rect 82967 53313 83045 53359
rect 83091 53313 83169 53359
rect 83215 53313 83293 53359
rect 83339 53313 83417 53359
rect 83463 53313 83541 53359
rect 83587 53313 83665 53359
rect 83711 53313 83789 53359
rect 83835 53313 83913 53359
rect 83959 53313 84037 53359
rect 84083 53313 84161 53359
rect 84207 53313 84285 53359
rect 84331 53313 84409 53359
rect 84455 53313 84533 53359
rect 84579 53313 84657 53359
rect 84703 53313 84781 53359
rect 84827 53313 84905 53359
rect 84951 53313 85029 53359
rect 85075 53313 85153 53359
rect 85199 53313 85277 53359
rect 85323 53313 85401 53359
rect 85447 53313 85525 53359
rect 85571 53313 85649 53359
rect 85695 53313 85706 53359
rect 0 53235 85706 53313
rect 0 53189 89 53235
rect 135 53189 213 53235
rect 259 53189 337 53235
rect 383 53189 461 53235
rect 507 53189 585 53235
rect 631 53189 709 53235
rect 755 53189 833 53235
rect 879 53189 957 53235
rect 1003 53189 1081 53235
rect 1127 53189 1205 53235
rect 1251 53189 1329 53235
rect 1375 53189 1453 53235
rect 1499 53189 1577 53235
rect 1623 53189 1701 53235
rect 1747 53189 1825 53235
rect 1871 53189 1949 53235
rect 1995 53189 2073 53235
rect 2119 53189 2197 53235
rect 2243 53189 2321 53235
rect 2367 53189 2445 53235
rect 2491 53189 2569 53235
rect 2615 53189 2693 53235
rect 2739 53189 2817 53235
rect 2863 53189 2941 53235
rect 2987 53189 3065 53235
rect 3111 53189 3189 53235
rect 3235 53189 3313 53235
rect 3359 53189 3437 53235
rect 3483 53189 3561 53235
rect 3607 53189 3685 53235
rect 3731 53189 3809 53235
rect 3855 53189 3933 53235
rect 3979 53189 4057 53235
rect 4103 53189 4181 53235
rect 4227 53189 4305 53235
rect 4351 53189 4429 53235
rect 4475 53189 4553 53235
rect 4599 53189 4677 53235
rect 4723 53189 4801 53235
rect 4847 53189 4925 53235
rect 4971 53189 5049 53235
rect 5095 53189 5173 53235
rect 5219 53189 5297 53235
rect 5343 53189 5421 53235
rect 5467 53189 5545 53235
rect 5591 53189 5669 53235
rect 5715 53189 5793 53235
rect 5839 53189 5917 53235
rect 5963 53189 6041 53235
rect 6087 53189 6165 53235
rect 6211 53189 6289 53235
rect 6335 53189 6413 53235
rect 6459 53189 6537 53235
rect 6583 53189 6661 53235
rect 6707 53189 6785 53235
rect 6831 53189 6909 53235
rect 6955 53189 7033 53235
rect 7079 53189 7157 53235
rect 7203 53189 7281 53235
rect 7327 53189 7405 53235
rect 7451 53189 7529 53235
rect 7575 53189 7653 53235
rect 7699 53189 7777 53235
rect 7823 53189 7901 53235
rect 7947 53189 8025 53235
rect 8071 53189 8149 53235
rect 8195 53189 8273 53235
rect 8319 53189 8397 53235
rect 8443 53189 8521 53235
rect 8567 53189 8645 53235
rect 8691 53189 8769 53235
rect 8815 53189 8893 53235
rect 8939 53189 9017 53235
rect 9063 53189 9141 53235
rect 9187 53189 9265 53235
rect 9311 53189 9389 53235
rect 9435 53189 9513 53235
rect 9559 53189 9637 53235
rect 9683 53189 9761 53235
rect 9807 53189 9885 53235
rect 9931 53189 10009 53235
rect 10055 53189 10133 53235
rect 10179 53189 10257 53235
rect 10303 53189 10381 53235
rect 10427 53189 10505 53235
rect 10551 53189 10629 53235
rect 10675 53189 10753 53235
rect 10799 53189 10877 53235
rect 10923 53189 11001 53235
rect 11047 53189 11125 53235
rect 11171 53189 11249 53235
rect 11295 53189 11373 53235
rect 11419 53189 11497 53235
rect 11543 53189 11621 53235
rect 11667 53189 11745 53235
rect 11791 53189 11869 53235
rect 11915 53189 11993 53235
rect 12039 53189 12117 53235
rect 12163 53189 12241 53235
rect 12287 53189 12365 53235
rect 12411 53189 12489 53235
rect 12535 53189 12613 53235
rect 12659 53189 12737 53235
rect 12783 53189 12861 53235
rect 12907 53189 12985 53235
rect 13031 53189 13109 53235
rect 13155 53189 13233 53235
rect 13279 53189 13357 53235
rect 13403 53189 13481 53235
rect 13527 53189 13605 53235
rect 13651 53189 13729 53235
rect 13775 53189 13853 53235
rect 13899 53189 13977 53235
rect 14023 53189 14101 53235
rect 14147 53189 14225 53235
rect 14271 53189 14349 53235
rect 14395 53189 14473 53235
rect 14519 53189 14597 53235
rect 14643 53189 14721 53235
rect 14767 53189 14845 53235
rect 14891 53189 14969 53235
rect 15015 53189 15093 53235
rect 15139 53189 15217 53235
rect 15263 53189 15341 53235
rect 15387 53189 15465 53235
rect 15511 53189 15589 53235
rect 15635 53189 15713 53235
rect 15759 53189 15837 53235
rect 15883 53189 15961 53235
rect 16007 53189 16085 53235
rect 16131 53189 16209 53235
rect 16255 53189 16333 53235
rect 16379 53189 16457 53235
rect 16503 53189 16581 53235
rect 16627 53189 16705 53235
rect 16751 53189 16829 53235
rect 16875 53189 16953 53235
rect 16999 53189 17077 53235
rect 17123 53189 17201 53235
rect 17247 53189 17325 53235
rect 17371 53189 17449 53235
rect 17495 53189 17573 53235
rect 17619 53189 17697 53235
rect 17743 53189 17821 53235
rect 17867 53189 17945 53235
rect 17991 53189 18069 53235
rect 18115 53189 18193 53235
rect 18239 53189 18317 53235
rect 18363 53189 18441 53235
rect 18487 53189 18565 53235
rect 18611 53189 18689 53235
rect 18735 53189 18813 53235
rect 18859 53189 18937 53235
rect 18983 53189 19061 53235
rect 19107 53189 19185 53235
rect 19231 53189 19309 53235
rect 19355 53189 19433 53235
rect 19479 53189 19557 53235
rect 19603 53189 19681 53235
rect 19727 53189 19805 53235
rect 19851 53189 19929 53235
rect 19975 53189 20053 53235
rect 20099 53189 20177 53235
rect 20223 53189 20301 53235
rect 20347 53189 20425 53235
rect 20471 53189 20549 53235
rect 20595 53189 20673 53235
rect 20719 53189 20797 53235
rect 20843 53189 20921 53235
rect 20967 53189 21045 53235
rect 21091 53189 21169 53235
rect 21215 53189 21293 53235
rect 21339 53189 21417 53235
rect 21463 53189 21541 53235
rect 21587 53189 21665 53235
rect 21711 53189 21789 53235
rect 21835 53189 21913 53235
rect 21959 53189 22037 53235
rect 22083 53189 22161 53235
rect 22207 53189 22285 53235
rect 22331 53189 22409 53235
rect 22455 53189 22533 53235
rect 22579 53189 22657 53235
rect 22703 53189 22781 53235
rect 22827 53189 22905 53235
rect 22951 53189 23029 53235
rect 23075 53189 23153 53235
rect 23199 53189 23277 53235
rect 23323 53189 23401 53235
rect 23447 53189 23525 53235
rect 23571 53189 23649 53235
rect 23695 53189 23773 53235
rect 23819 53189 23897 53235
rect 23943 53189 24021 53235
rect 24067 53189 24145 53235
rect 24191 53189 24269 53235
rect 24315 53189 24393 53235
rect 24439 53189 24517 53235
rect 24563 53189 24641 53235
rect 24687 53189 24765 53235
rect 24811 53189 24889 53235
rect 24935 53189 25013 53235
rect 25059 53189 25137 53235
rect 25183 53189 25261 53235
rect 25307 53189 25385 53235
rect 25431 53189 25509 53235
rect 25555 53189 25633 53235
rect 25679 53189 25757 53235
rect 25803 53189 25881 53235
rect 25927 53189 26005 53235
rect 26051 53189 26129 53235
rect 26175 53189 26253 53235
rect 26299 53189 26377 53235
rect 26423 53189 26501 53235
rect 26547 53189 26625 53235
rect 26671 53189 26749 53235
rect 26795 53189 26873 53235
rect 26919 53189 26997 53235
rect 27043 53189 27121 53235
rect 27167 53189 27245 53235
rect 27291 53189 27369 53235
rect 27415 53189 27493 53235
rect 27539 53189 27617 53235
rect 27663 53189 27741 53235
rect 27787 53189 27865 53235
rect 27911 53189 27989 53235
rect 28035 53189 28113 53235
rect 28159 53189 28237 53235
rect 28283 53189 28361 53235
rect 28407 53189 28485 53235
rect 28531 53189 28609 53235
rect 28655 53189 28733 53235
rect 28779 53189 28857 53235
rect 28903 53189 28981 53235
rect 29027 53189 29105 53235
rect 29151 53189 29229 53235
rect 29275 53189 29353 53235
rect 29399 53189 29477 53235
rect 29523 53189 29601 53235
rect 29647 53189 29725 53235
rect 29771 53189 29849 53235
rect 29895 53189 29973 53235
rect 30019 53189 30097 53235
rect 30143 53189 30221 53235
rect 30267 53189 30345 53235
rect 30391 53189 30469 53235
rect 30515 53189 30593 53235
rect 30639 53189 30717 53235
rect 30763 53189 30841 53235
rect 30887 53189 30965 53235
rect 31011 53189 31089 53235
rect 31135 53189 31213 53235
rect 31259 53189 31337 53235
rect 31383 53189 31461 53235
rect 31507 53189 31585 53235
rect 31631 53189 31709 53235
rect 31755 53189 31833 53235
rect 31879 53189 31957 53235
rect 32003 53189 32081 53235
rect 32127 53189 32205 53235
rect 32251 53189 32329 53235
rect 32375 53189 32453 53235
rect 32499 53189 32577 53235
rect 32623 53189 32701 53235
rect 32747 53189 32825 53235
rect 32871 53189 32949 53235
rect 32995 53189 33073 53235
rect 33119 53189 33197 53235
rect 33243 53189 33321 53235
rect 33367 53189 33445 53235
rect 33491 53189 33569 53235
rect 33615 53189 33693 53235
rect 33739 53189 33817 53235
rect 33863 53189 33941 53235
rect 33987 53189 34065 53235
rect 34111 53189 34189 53235
rect 34235 53189 34313 53235
rect 34359 53189 34437 53235
rect 34483 53189 34561 53235
rect 34607 53189 34685 53235
rect 34731 53189 34809 53235
rect 34855 53189 34933 53235
rect 34979 53189 35057 53235
rect 35103 53189 35181 53235
rect 35227 53189 35305 53235
rect 35351 53189 35429 53235
rect 35475 53189 35553 53235
rect 35599 53189 35677 53235
rect 35723 53189 35801 53235
rect 35847 53189 35925 53235
rect 35971 53189 36049 53235
rect 36095 53189 36173 53235
rect 36219 53189 36297 53235
rect 36343 53189 36421 53235
rect 36467 53189 36545 53235
rect 36591 53189 36669 53235
rect 36715 53189 36793 53235
rect 36839 53189 36917 53235
rect 36963 53189 37041 53235
rect 37087 53189 37165 53235
rect 37211 53189 37289 53235
rect 37335 53189 37413 53235
rect 37459 53189 37537 53235
rect 37583 53189 37661 53235
rect 37707 53189 37785 53235
rect 37831 53189 37909 53235
rect 37955 53189 38033 53235
rect 38079 53189 38157 53235
rect 38203 53189 38281 53235
rect 38327 53189 38405 53235
rect 38451 53189 38529 53235
rect 38575 53189 38653 53235
rect 38699 53189 38777 53235
rect 38823 53189 38901 53235
rect 38947 53189 39025 53235
rect 39071 53189 39149 53235
rect 39195 53189 39273 53235
rect 39319 53189 39397 53235
rect 39443 53189 39521 53235
rect 39567 53189 39645 53235
rect 39691 53189 39769 53235
rect 39815 53189 39893 53235
rect 39939 53189 40017 53235
rect 40063 53189 40141 53235
rect 40187 53189 40265 53235
rect 40311 53189 40389 53235
rect 40435 53189 40513 53235
rect 40559 53189 40637 53235
rect 40683 53189 40761 53235
rect 40807 53189 40885 53235
rect 40931 53189 41009 53235
rect 41055 53189 41133 53235
rect 41179 53189 41257 53235
rect 41303 53189 41381 53235
rect 41427 53189 41505 53235
rect 41551 53189 41629 53235
rect 41675 53189 41753 53235
rect 41799 53189 41877 53235
rect 41923 53189 42001 53235
rect 42047 53189 42125 53235
rect 42171 53189 42249 53235
rect 42295 53189 42373 53235
rect 42419 53189 42497 53235
rect 42543 53189 42621 53235
rect 42667 53189 42745 53235
rect 42791 53189 42869 53235
rect 42915 53189 42993 53235
rect 43039 53189 43117 53235
rect 43163 53189 43241 53235
rect 43287 53189 43365 53235
rect 43411 53189 43489 53235
rect 43535 53189 43613 53235
rect 43659 53189 43737 53235
rect 43783 53189 43861 53235
rect 43907 53189 43985 53235
rect 44031 53189 44109 53235
rect 44155 53189 44233 53235
rect 44279 53189 44357 53235
rect 44403 53189 44481 53235
rect 44527 53189 44605 53235
rect 44651 53189 44729 53235
rect 44775 53189 44853 53235
rect 44899 53189 44977 53235
rect 45023 53189 45101 53235
rect 45147 53189 45225 53235
rect 45271 53189 45349 53235
rect 45395 53189 45473 53235
rect 45519 53189 45597 53235
rect 45643 53189 45721 53235
rect 45767 53189 45845 53235
rect 45891 53189 45969 53235
rect 46015 53189 46093 53235
rect 46139 53189 46217 53235
rect 46263 53189 46341 53235
rect 46387 53189 46465 53235
rect 46511 53189 46589 53235
rect 46635 53189 46713 53235
rect 46759 53189 46837 53235
rect 46883 53189 46961 53235
rect 47007 53189 47085 53235
rect 47131 53189 47209 53235
rect 47255 53189 47333 53235
rect 47379 53189 47457 53235
rect 47503 53189 47581 53235
rect 47627 53189 47705 53235
rect 47751 53189 47829 53235
rect 47875 53189 47953 53235
rect 47999 53189 48077 53235
rect 48123 53189 48201 53235
rect 48247 53189 48325 53235
rect 48371 53189 48449 53235
rect 48495 53189 48573 53235
rect 48619 53189 48697 53235
rect 48743 53189 48821 53235
rect 48867 53189 48945 53235
rect 48991 53189 49069 53235
rect 49115 53189 49193 53235
rect 49239 53189 49317 53235
rect 49363 53189 49441 53235
rect 49487 53189 49565 53235
rect 49611 53189 49689 53235
rect 49735 53189 49813 53235
rect 49859 53189 49937 53235
rect 49983 53189 50061 53235
rect 50107 53189 50185 53235
rect 50231 53189 50309 53235
rect 50355 53189 50433 53235
rect 50479 53189 50557 53235
rect 50603 53189 50681 53235
rect 50727 53189 50805 53235
rect 50851 53189 50929 53235
rect 50975 53189 51053 53235
rect 51099 53189 51177 53235
rect 51223 53189 51301 53235
rect 51347 53189 51425 53235
rect 51471 53189 51549 53235
rect 51595 53189 51673 53235
rect 51719 53189 51797 53235
rect 51843 53189 51921 53235
rect 51967 53189 52045 53235
rect 52091 53189 52169 53235
rect 52215 53189 52293 53235
rect 52339 53189 52417 53235
rect 52463 53189 52541 53235
rect 52587 53189 52665 53235
rect 52711 53189 52789 53235
rect 52835 53189 52913 53235
rect 52959 53189 53037 53235
rect 53083 53189 53161 53235
rect 53207 53189 53285 53235
rect 53331 53189 53409 53235
rect 53455 53189 53533 53235
rect 53579 53189 53657 53235
rect 53703 53189 53781 53235
rect 53827 53189 53905 53235
rect 53951 53189 54029 53235
rect 54075 53189 54153 53235
rect 54199 53189 54277 53235
rect 54323 53189 54401 53235
rect 54447 53189 54525 53235
rect 54571 53189 54649 53235
rect 54695 53189 54773 53235
rect 54819 53189 54897 53235
rect 54943 53189 55021 53235
rect 55067 53189 55145 53235
rect 55191 53189 55269 53235
rect 55315 53189 55393 53235
rect 55439 53189 55517 53235
rect 55563 53189 55641 53235
rect 55687 53189 55765 53235
rect 55811 53189 55889 53235
rect 55935 53189 56013 53235
rect 56059 53189 56137 53235
rect 56183 53189 56261 53235
rect 56307 53189 56385 53235
rect 56431 53189 56509 53235
rect 56555 53189 56633 53235
rect 56679 53189 56757 53235
rect 56803 53189 56881 53235
rect 56927 53189 57005 53235
rect 57051 53189 57129 53235
rect 57175 53189 57253 53235
rect 57299 53189 57377 53235
rect 57423 53189 57501 53235
rect 57547 53189 57625 53235
rect 57671 53189 57749 53235
rect 57795 53189 57873 53235
rect 57919 53189 57997 53235
rect 58043 53189 58121 53235
rect 58167 53189 58245 53235
rect 58291 53189 58369 53235
rect 58415 53189 58493 53235
rect 58539 53189 58617 53235
rect 58663 53189 58741 53235
rect 58787 53189 58865 53235
rect 58911 53189 58989 53235
rect 59035 53189 59113 53235
rect 59159 53189 59237 53235
rect 59283 53189 59361 53235
rect 59407 53189 59485 53235
rect 59531 53189 59609 53235
rect 59655 53189 59733 53235
rect 59779 53189 59857 53235
rect 59903 53189 59981 53235
rect 60027 53189 60105 53235
rect 60151 53189 60229 53235
rect 60275 53189 60353 53235
rect 60399 53189 60477 53235
rect 60523 53189 60601 53235
rect 60647 53189 60725 53235
rect 60771 53189 60849 53235
rect 60895 53189 60973 53235
rect 61019 53189 61097 53235
rect 61143 53189 61221 53235
rect 61267 53189 61345 53235
rect 61391 53189 61469 53235
rect 61515 53189 61593 53235
rect 61639 53189 61717 53235
rect 61763 53189 61841 53235
rect 61887 53189 61965 53235
rect 62011 53189 62089 53235
rect 62135 53189 62213 53235
rect 62259 53189 62337 53235
rect 62383 53189 62461 53235
rect 62507 53189 62585 53235
rect 62631 53189 62709 53235
rect 62755 53189 62833 53235
rect 62879 53189 62957 53235
rect 63003 53189 63081 53235
rect 63127 53189 63205 53235
rect 63251 53189 63329 53235
rect 63375 53189 63453 53235
rect 63499 53189 63577 53235
rect 63623 53189 63701 53235
rect 63747 53189 63825 53235
rect 63871 53189 63949 53235
rect 63995 53189 64073 53235
rect 64119 53189 64197 53235
rect 64243 53189 64321 53235
rect 64367 53189 64445 53235
rect 64491 53189 64569 53235
rect 64615 53189 64693 53235
rect 64739 53189 64817 53235
rect 64863 53189 64941 53235
rect 64987 53189 65065 53235
rect 65111 53189 65189 53235
rect 65235 53189 65313 53235
rect 65359 53189 65437 53235
rect 65483 53189 65561 53235
rect 65607 53189 65685 53235
rect 65731 53189 65809 53235
rect 65855 53189 65933 53235
rect 65979 53189 66057 53235
rect 66103 53189 66181 53235
rect 66227 53189 66305 53235
rect 66351 53189 66429 53235
rect 66475 53189 66553 53235
rect 66599 53189 66677 53235
rect 66723 53189 66801 53235
rect 66847 53189 66925 53235
rect 66971 53189 67049 53235
rect 67095 53189 67173 53235
rect 67219 53189 67297 53235
rect 67343 53189 67421 53235
rect 67467 53189 67545 53235
rect 67591 53189 67669 53235
rect 67715 53189 67793 53235
rect 67839 53189 67917 53235
rect 67963 53189 68041 53235
rect 68087 53189 68165 53235
rect 68211 53189 68289 53235
rect 68335 53189 68413 53235
rect 68459 53189 68537 53235
rect 68583 53189 68661 53235
rect 68707 53189 68785 53235
rect 68831 53189 68909 53235
rect 68955 53189 69033 53235
rect 69079 53189 69157 53235
rect 69203 53189 69281 53235
rect 69327 53189 69405 53235
rect 69451 53189 69529 53235
rect 69575 53189 69653 53235
rect 69699 53189 69777 53235
rect 69823 53189 69901 53235
rect 69947 53189 70025 53235
rect 70071 53189 70149 53235
rect 70195 53189 70273 53235
rect 70319 53189 70397 53235
rect 70443 53189 70521 53235
rect 70567 53189 70645 53235
rect 70691 53189 70769 53235
rect 70815 53189 70893 53235
rect 70939 53189 71017 53235
rect 71063 53189 71141 53235
rect 71187 53189 71265 53235
rect 71311 53189 71389 53235
rect 71435 53189 71513 53235
rect 71559 53189 71637 53235
rect 71683 53189 71761 53235
rect 71807 53189 71885 53235
rect 71931 53189 72009 53235
rect 72055 53189 72133 53235
rect 72179 53189 72257 53235
rect 72303 53189 72381 53235
rect 72427 53189 72505 53235
rect 72551 53189 72629 53235
rect 72675 53189 72753 53235
rect 72799 53189 72877 53235
rect 72923 53189 73001 53235
rect 73047 53189 73125 53235
rect 73171 53189 73249 53235
rect 73295 53189 73373 53235
rect 73419 53189 73497 53235
rect 73543 53189 73621 53235
rect 73667 53189 73745 53235
rect 73791 53189 73869 53235
rect 73915 53189 73993 53235
rect 74039 53189 74117 53235
rect 74163 53189 74241 53235
rect 74287 53189 74365 53235
rect 74411 53189 74489 53235
rect 74535 53189 74613 53235
rect 74659 53189 74737 53235
rect 74783 53189 74861 53235
rect 74907 53189 74985 53235
rect 75031 53189 75109 53235
rect 75155 53189 75233 53235
rect 75279 53189 75357 53235
rect 75403 53189 75481 53235
rect 75527 53189 75605 53235
rect 75651 53189 75729 53235
rect 75775 53189 75853 53235
rect 75899 53189 75977 53235
rect 76023 53189 76101 53235
rect 76147 53189 76225 53235
rect 76271 53189 76349 53235
rect 76395 53189 76473 53235
rect 76519 53189 76597 53235
rect 76643 53189 76721 53235
rect 76767 53189 76845 53235
rect 76891 53189 76969 53235
rect 77015 53189 77093 53235
rect 77139 53189 77217 53235
rect 77263 53189 77341 53235
rect 77387 53189 77465 53235
rect 77511 53189 77589 53235
rect 77635 53189 77713 53235
rect 77759 53189 77837 53235
rect 77883 53189 77961 53235
rect 78007 53189 78085 53235
rect 78131 53189 78209 53235
rect 78255 53189 78333 53235
rect 78379 53189 78457 53235
rect 78503 53189 78581 53235
rect 78627 53189 78705 53235
rect 78751 53189 78829 53235
rect 78875 53189 78953 53235
rect 78999 53189 79077 53235
rect 79123 53189 79201 53235
rect 79247 53189 79325 53235
rect 79371 53189 79449 53235
rect 79495 53189 79573 53235
rect 79619 53189 79697 53235
rect 79743 53189 79821 53235
rect 79867 53189 79945 53235
rect 79991 53189 80069 53235
rect 80115 53189 80193 53235
rect 80239 53189 80317 53235
rect 80363 53189 80441 53235
rect 80487 53189 80565 53235
rect 80611 53189 80689 53235
rect 80735 53189 80813 53235
rect 80859 53189 80937 53235
rect 80983 53189 81061 53235
rect 81107 53189 81185 53235
rect 81231 53189 81309 53235
rect 81355 53189 81433 53235
rect 81479 53189 81557 53235
rect 81603 53189 81681 53235
rect 81727 53189 81805 53235
rect 81851 53189 81929 53235
rect 81975 53189 82053 53235
rect 82099 53189 82177 53235
rect 82223 53189 82301 53235
rect 82347 53189 82425 53235
rect 82471 53189 82549 53235
rect 82595 53189 82673 53235
rect 82719 53189 82797 53235
rect 82843 53189 82921 53235
rect 82967 53189 83045 53235
rect 83091 53189 83169 53235
rect 83215 53189 83293 53235
rect 83339 53189 83417 53235
rect 83463 53189 83541 53235
rect 83587 53189 83665 53235
rect 83711 53189 83789 53235
rect 83835 53189 83913 53235
rect 83959 53189 84037 53235
rect 84083 53189 84161 53235
rect 84207 53189 84285 53235
rect 84331 53189 84409 53235
rect 84455 53189 84533 53235
rect 84579 53189 84657 53235
rect 84703 53189 84781 53235
rect 84827 53189 84905 53235
rect 84951 53189 85029 53235
rect 85075 53189 85153 53235
rect 85199 53189 85277 53235
rect 85323 53189 85401 53235
rect 85447 53189 85525 53235
rect 85571 53189 85649 53235
rect 85695 53189 85706 53235
rect 0 53111 85706 53189
rect 0 53065 89 53111
rect 135 53065 213 53111
rect 259 53065 337 53111
rect 383 53065 461 53111
rect 507 53065 585 53111
rect 631 53065 709 53111
rect 755 53065 833 53111
rect 879 53065 957 53111
rect 1003 53065 1081 53111
rect 1127 53065 1205 53111
rect 1251 53065 1329 53111
rect 1375 53065 1453 53111
rect 1499 53065 1577 53111
rect 1623 53065 1701 53111
rect 1747 53065 1825 53111
rect 1871 53065 1949 53111
rect 1995 53065 2073 53111
rect 2119 53065 2197 53111
rect 2243 53065 2321 53111
rect 2367 53065 2445 53111
rect 2491 53065 2569 53111
rect 2615 53065 2693 53111
rect 2739 53065 2817 53111
rect 2863 53065 2941 53111
rect 2987 53065 3065 53111
rect 3111 53065 3189 53111
rect 3235 53065 3313 53111
rect 3359 53065 3437 53111
rect 3483 53065 3561 53111
rect 3607 53065 3685 53111
rect 3731 53065 3809 53111
rect 3855 53065 3933 53111
rect 3979 53065 4057 53111
rect 4103 53065 4181 53111
rect 4227 53065 4305 53111
rect 4351 53065 4429 53111
rect 4475 53065 4553 53111
rect 4599 53065 4677 53111
rect 4723 53065 4801 53111
rect 4847 53065 4925 53111
rect 4971 53065 5049 53111
rect 5095 53065 5173 53111
rect 5219 53065 5297 53111
rect 5343 53065 5421 53111
rect 5467 53065 5545 53111
rect 5591 53065 5669 53111
rect 5715 53065 5793 53111
rect 5839 53065 5917 53111
rect 5963 53065 6041 53111
rect 6087 53065 6165 53111
rect 6211 53065 6289 53111
rect 6335 53065 6413 53111
rect 6459 53065 6537 53111
rect 6583 53065 6661 53111
rect 6707 53065 6785 53111
rect 6831 53065 6909 53111
rect 6955 53065 7033 53111
rect 7079 53065 7157 53111
rect 7203 53065 7281 53111
rect 7327 53065 7405 53111
rect 7451 53065 7529 53111
rect 7575 53065 7653 53111
rect 7699 53065 7777 53111
rect 7823 53065 7901 53111
rect 7947 53065 8025 53111
rect 8071 53065 8149 53111
rect 8195 53065 8273 53111
rect 8319 53065 8397 53111
rect 8443 53065 8521 53111
rect 8567 53065 8645 53111
rect 8691 53065 8769 53111
rect 8815 53065 8893 53111
rect 8939 53065 9017 53111
rect 9063 53065 9141 53111
rect 9187 53065 9265 53111
rect 9311 53065 9389 53111
rect 9435 53065 9513 53111
rect 9559 53065 9637 53111
rect 9683 53065 9761 53111
rect 9807 53065 9885 53111
rect 9931 53065 10009 53111
rect 10055 53065 10133 53111
rect 10179 53065 10257 53111
rect 10303 53065 10381 53111
rect 10427 53065 10505 53111
rect 10551 53065 10629 53111
rect 10675 53065 10753 53111
rect 10799 53065 10877 53111
rect 10923 53065 11001 53111
rect 11047 53065 11125 53111
rect 11171 53065 11249 53111
rect 11295 53065 11373 53111
rect 11419 53065 11497 53111
rect 11543 53065 11621 53111
rect 11667 53065 11745 53111
rect 11791 53065 11869 53111
rect 11915 53065 11993 53111
rect 12039 53065 12117 53111
rect 12163 53065 12241 53111
rect 12287 53065 12365 53111
rect 12411 53065 12489 53111
rect 12535 53065 12613 53111
rect 12659 53065 12737 53111
rect 12783 53065 12861 53111
rect 12907 53065 12985 53111
rect 13031 53065 13109 53111
rect 13155 53065 13233 53111
rect 13279 53065 13357 53111
rect 13403 53065 13481 53111
rect 13527 53065 13605 53111
rect 13651 53065 13729 53111
rect 13775 53065 13853 53111
rect 13899 53065 13977 53111
rect 14023 53065 14101 53111
rect 14147 53065 14225 53111
rect 14271 53065 14349 53111
rect 14395 53065 14473 53111
rect 14519 53065 14597 53111
rect 14643 53065 14721 53111
rect 14767 53065 14845 53111
rect 14891 53065 14969 53111
rect 15015 53065 15093 53111
rect 15139 53065 15217 53111
rect 15263 53065 15341 53111
rect 15387 53065 15465 53111
rect 15511 53065 15589 53111
rect 15635 53065 15713 53111
rect 15759 53065 15837 53111
rect 15883 53065 15961 53111
rect 16007 53065 16085 53111
rect 16131 53065 16209 53111
rect 16255 53065 16333 53111
rect 16379 53065 16457 53111
rect 16503 53065 16581 53111
rect 16627 53065 16705 53111
rect 16751 53065 16829 53111
rect 16875 53065 16953 53111
rect 16999 53065 17077 53111
rect 17123 53065 17201 53111
rect 17247 53065 17325 53111
rect 17371 53065 17449 53111
rect 17495 53065 17573 53111
rect 17619 53065 17697 53111
rect 17743 53065 17821 53111
rect 17867 53065 17945 53111
rect 17991 53065 18069 53111
rect 18115 53065 18193 53111
rect 18239 53065 18317 53111
rect 18363 53065 18441 53111
rect 18487 53065 18565 53111
rect 18611 53065 18689 53111
rect 18735 53065 18813 53111
rect 18859 53065 18937 53111
rect 18983 53065 19061 53111
rect 19107 53065 19185 53111
rect 19231 53065 19309 53111
rect 19355 53065 19433 53111
rect 19479 53065 19557 53111
rect 19603 53065 19681 53111
rect 19727 53065 19805 53111
rect 19851 53065 19929 53111
rect 19975 53065 20053 53111
rect 20099 53065 20177 53111
rect 20223 53065 20301 53111
rect 20347 53065 20425 53111
rect 20471 53065 20549 53111
rect 20595 53065 20673 53111
rect 20719 53065 20797 53111
rect 20843 53065 20921 53111
rect 20967 53065 21045 53111
rect 21091 53065 21169 53111
rect 21215 53065 21293 53111
rect 21339 53065 21417 53111
rect 21463 53065 21541 53111
rect 21587 53065 21665 53111
rect 21711 53065 21789 53111
rect 21835 53065 21913 53111
rect 21959 53065 22037 53111
rect 22083 53065 22161 53111
rect 22207 53065 22285 53111
rect 22331 53065 22409 53111
rect 22455 53065 22533 53111
rect 22579 53065 22657 53111
rect 22703 53065 22781 53111
rect 22827 53065 22905 53111
rect 22951 53065 23029 53111
rect 23075 53065 23153 53111
rect 23199 53065 23277 53111
rect 23323 53065 23401 53111
rect 23447 53065 23525 53111
rect 23571 53065 23649 53111
rect 23695 53065 23773 53111
rect 23819 53065 23897 53111
rect 23943 53065 24021 53111
rect 24067 53065 24145 53111
rect 24191 53065 24269 53111
rect 24315 53065 24393 53111
rect 24439 53065 24517 53111
rect 24563 53065 24641 53111
rect 24687 53065 24765 53111
rect 24811 53065 24889 53111
rect 24935 53065 25013 53111
rect 25059 53065 25137 53111
rect 25183 53065 25261 53111
rect 25307 53065 25385 53111
rect 25431 53065 25509 53111
rect 25555 53065 25633 53111
rect 25679 53065 25757 53111
rect 25803 53065 25881 53111
rect 25927 53065 26005 53111
rect 26051 53065 26129 53111
rect 26175 53065 26253 53111
rect 26299 53065 26377 53111
rect 26423 53065 26501 53111
rect 26547 53065 26625 53111
rect 26671 53065 26749 53111
rect 26795 53065 26873 53111
rect 26919 53065 26997 53111
rect 27043 53065 27121 53111
rect 27167 53065 27245 53111
rect 27291 53065 27369 53111
rect 27415 53065 27493 53111
rect 27539 53065 27617 53111
rect 27663 53065 27741 53111
rect 27787 53065 27865 53111
rect 27911 53065 27989 53111
rect 28035 53065 28113 53111
rect 28159 53065 28237 53111
rect 28283 53065 28361 53111
rect 28407 53065 28485 53111
rect 28531 53065 28609 53111
rect 28655 53065 28733 53111
rect 28779 53065 28857 53111
rect 28903 53065 28981 53111
rect 29027 53065 29105 53111
rect 29151 53065 29229 53111
rect 29275 53065 29353 53111
rect 29399 53065 29477 53111
rect 29523 53065 29601 53111
rect 29647 53065 29725 53111
rect 29771 53065 29849 53111
rect 29895 53065 29973 53111
rect 30019 53065 30097 53111
rect 30143 53065 30221 53111
rect 30267 53065 30345 53111
rect 30391 53065 30469 53111
rect 30515 53065 30593 53111
rect 30639 53065 30717 53111
rect 30763 53065 30841 53111
rect 30887 53065 30965 53111
rect 31011 53065 31089 53111
rect 31135 53065 31213 53111
rect 31259 53065 31337 53111
rect 31383 53065 31461 53111
rect 31507 53065 31585 53111
rect 31631 53065 31709 53111
rect 31755 53065 31833 53111
rect 31879 53065 31957 53111
rect 32003 53065 32081 53111
rect 32127 53065 32205 53111
rect 32251 53065 32329 53111
rect 32375 53065 32453 53111
rect 32499 53065 32577 53111
rect 32623 53065 32701 53111
rect 32747 53065 32825 53111
rect 32871 53065 32949 53111
rect 32995 53065 33073 53111
rect 33119 53065 33197 53111
rect 33243 53065 33321 53111
rect 33367 53065 33445 53111
rect 33491 53065 33569 53111
rect 33615 53065 33693 53111
rect 33739 53065 33817 53111
rect 33863 53065 33941 53111
rect 33987 53065 34065 53111
rect 34111 53065 34189 53111
rect 34235 53065 34313 53111
rect 34359 53065 34437 53111
rect 34483 53065 34561 53111
rect 34607 53065 34685 53111
rect 34731 53065 34809 53111
rect 34855 53065 34933 53111
rect 34979 53065 35057 53111
rect 35103 53065 35181 53111
rect 35227 53065 35305 53111
rect 35351 53065 35429 53111
rect 35475 53065 35553 53111
rect 35599 53065 35677 53111
rect 35723 53065 35801 53111
rect 35847 53065 35925 53111
rect 35971 53065 36049 53111
rect 36095 53065 36173 53111
rect 36219 53065 36297 53111
rect 36343 53065 36421 53111
rect 36467 53065 36545 53111
rect 36591 53065 36669 53111
rect 36715 53065 36793 53111
rect 36839 53065 36917 53111
rect 36963 53065 37041 53111
rect 37087 53065 37165 53111
rect 37211 53065 37289 53111
rect 37335 53065 37413 53111
rect 37459 53065 37537 53111
rect 37583 53065 37661 53111
rect 37707 53065 37785 53111
rect 37831 53065 37909 53111
rect 37955 53065 38033 53111
rect 38079 53065 38157 53111
rect 38203 53065 38281 53111
rect 38327 53065 38405 53111
rect 38451 53065 38529 53111
rect 38575 53065 38653 53111
rect 38699 53065 38777 53111
rect 38823 53065 38901 53111
rect 38947 53065 39025 53111
rect 39071 53065 39149 53111
rect 39195 53065 39273 53111
rect 39319 53065 39397 53111
rect 39443 53065 39521 53111
rect 39567 53065 39645 53111
rect 39691 53065 39769 53111
rect 39815 53065 39893 53111
rect 39939 53065 40017 53111
rect 40063 53065 40141 53111
rect 40187 53065 40265 53111
rect 40311 53065 40389 53111
rect 40435 53065 40513 53111
rect 40559 53065 40637 53111
rect 40683 53065 40761 53111
rect 40807 53065 40885 53111
rect 40931 53065 41009 53111
rect 41055 53065 41133 53111
rect 41179 53065 41257 53111
rect 41303 53065 41381 53111
rect 41427 53065 41505 53111
rect 41551 53065 41629 53111
rect 41675 53065 41753 53111
rect 41799 53065 41877 53111
rect 41923 53065 42001 53111
rect 42047 53065 42125 53111
rect 42171 53065 42249 53111
rect 42295 53065 42373 53111
rect 42419 53065 42497 53111
rect 42543 53065 42621 53111
rect 42667 53065 42745 53111
rect 42791 53065 42869 53111
rect 42915 53065 42993 53111
rect 43039 53065 43117 53111
rect 43163 53065 43241 53111
rect 43287 53065 43365 53111
rect 43411 53065 43489 53111
rect 43535 53065 43613 53111
rect 43659 53065 43737 53111
rect 43783 53065 43861 53111
rect 43907 53065 43985 53111
rect 44031 53065 44109 53111
rect 44155 53065 44233 53111
rect 44279 53065 44357 53111
rect 44403 53065 44481 53111
rect 44527 53065 44605 53111
rect 44651 53065 44729 53111
rect 44775 53065 44853 53111
rect 44899 53065 44977 53111
rect 45023 53065 45101 53111
rect 45147 53065 45225 53111
rect 45271 53065 45349 53111
rect 45395 53065 45473 53111
rect 45519 53065 45597 53111
rect 45643 53065 45721 53111
rect 45767 53065 45845 53111
rect 45891 53065 45969 53111
rect 46015 53065 46093 53111
rect 46139 53065 46217 53111
rect 46263 53065 46341 53111
rect 46387 53065 46465 53111
rect 46511 53065 46589 53111
rect 46635 53065 46713 53111
rect 46759 53065 46837 53111
rect 46883 53065 46961 53111
rect 47007 53065 47085 53111
rect 47131 53065 47209 53111
rect 47255 53065 47333 53111
rect 47379 53065 47457 53111
rect 47503 53065 47581 53111
rect 47627 53065 47705 53111
rect 47751 53065 47829 53111
rect 47875 53065 47953 53111
rect 47999 53065 48077 53111
rect 48123 53065 48201 53111
rect 48247 53065 48325 53111
rect 48371 53065 48449 53111
rect 48495 53065 48573 53111
rect 48619 53065 48697 53111
rect 48743 53065 48821 53111
rect 48867 53065 48945 53111
rect 48991 53065 49069 53111
rect 49115 53065 49193 53111
rect 49239 53065 49317 53111
rect 49363 53065 49441 53111
rect 49487 53065 49565 53111
rect 49611 53065 49689 53111
rect 49735 53065 49813 53111
rect 49859 53065 49937 53111
rect 49983 53065 50061 53111
rect 50107 53065 50185 53111
rect 50231 53065 50309 53111
rect 50355 53065 50433 53111
rect 50479 53065 50557 53111
rect 50603 53065 50681 53111
rect 50727 53065 50805 53111
rect 50851 53065 50929 53111
rect 50975 53065 51053 53111
rect 51099 53065 51177 53111
rect 51223 53065 51301 53111
rect 51347 53065 51425 53111
rect 51471 53065 51549 53111
rect 51595 53065 51673 53111
rect 51719 53065 51797 53111
rect 51843 53065 51921 53111
rect 51967 53065 52045 53111
rect 52091 53065 52169 53111
rect 52215 53065 52293 53111
rect 52339 53065 52417 53111
rect 52463 53065 52541 53111
rect 52587 53065 52665 53111
rect 52711 53065 52789 53111
rect 52835 53065 52913 53111
rect 52959 53065 53037 53111
rect 53083 53065 53161 53111
rect 53207 53065 53285 53111
rect 53331 53065 53409 53111
rect 53455 53065 53533 53111
rect 53579 53065 53657 53111
rect 53703 53065 53781 53111
rect 53827 53065 53905 53111
rect 53951 53065 54029 53111
rect 54075 53065 54153 53111
rect 54199 53065 54277 53111
rect 54323 53065 54401 53111
rect 54447 53065 54525 53111
rect 54571 53065 54649 53111
rect 54695 53065 54773 53111
rect 54819 53065 54897 53111
rect 54943 53065 55021 53111
rect 55067 53065 55145 53111
rect 55191 53065 55269 53111
rect 55315 53065 55393 53111
rect 55439 53065 55517 53111
rect 55563 53065 55641 53111
rect 55687 53065 55765 53111
rect 55811 53065 55889 53111
rect 55935 53065 56013 53111
rect 56059 53065 56137 53111
rect 56183 53065 56261 53111
rect 56307 53065 56385 53111
rect 56431 53065 56509 53111
rect 56555 53065 56633 53111
rect 56679 53065 56757 53111
rect 56803 53065 56881 53111
rect 56927 53065 57005 53111
rect 57051 53065 57129 53111
rect 57175 53065 57253 53111
rect 57299 53065 57377 53111
rect 57423 53065 57501 53111
rect 57547 53065 57625 53111
rect 57671 53065 57749 53111
rect 57795 53065 57873 53111
rect 57919 53065 57997 53111
rect 58043 53065 58121 53111
rect 58167 53065 58245 53111
rect 58291 53065 58369 53111
rect 58415 53065 58493 53111
rect 58539 53065 58617 53111
rect 58663 53065 58741 53111
rect 58787 53065 58865 53111
rect 58911 53065 58989 53111
rect 59035 53065 59113 53111
rect 59159 53065 59237 53111
rect 59283 53065 59361 53111
rect 59407 53065 59485 53111
rect 59531 53065 59609 53111
rect 59655 53065 59733 53111
rect 59779 53065 59857 53111
rect 59903 53065 59981 53111
rect 60027 53065 60105 53111
rect 60151 53065 60229 53111
rect 60275 53065 60353 53111
rect 60399 53065 60477 53111
rect 60523 53065 60601 53111
rect 60647 53065 60725 53111
rect 60771 53065 60849 53111
rect 60895 53065 60973 53111
rect 61019 53065 61097 53111
rect 61143 53065 61221 53111
rect 61267 53065 61345 53111
rect 61391 53065 61469 53111
rect 61515 53065 61593 53111
rect 61639 53065 61717 53111
rect 61763 53065 61841 53111
rect 61887 53065 61965 53111
rect 62011 53065 62089 53111
rect 62135 53065 62213 53111
rect 62259 53065 62337 53111
rect 62383 53065 62461 53111
rect 62507 53065 62585 53111
rect 62631 53065 62709 53111
rect 62755 53065 62833 53111
rect 62879 53065 62957 53111
rect 63003 53065 63081 53111
rect 63127 53065 63205 53111
rect 63251 53065 63329 53111
rect 63375 53065 63453 53111
rect 63499 53065 63577 53111
rect 63623 53065 63701 53111
rect 63747 53065 63825 53111
rect 63871 53065 63949 53111
rect 63995 53065 64073 53111
rect 64119 53065 64197 53111
rect 64243 53065 64321 53111
rect 64367 53065 64445 53111
rect 64491 53065 64569 53111
rect 64615 53065 64693 53111
rect 64739 53065 64817 53111
rect 64863 53065 64941 53111
rect 64987 53065 65065 53111
rect 65111 53065 65189 53111
rect 65235 53065 65313 53111
rect 65359 53065 65437 53111
rect 65483 53065 65561 53111
rect 65607 53065 65685 53111
rect 65731 53065 65809 53111
rect 65855 53065 65933 53111
rect 65979 53065 66057 53111
rect 66103 53065 66181 53111
rect 66227 53065 66305 53111
rect 66351 53065 66429 53111
rect 66475 53065 66553 53111
rect 66599 53065 66677 53111
rect 66723 53065 66801 53111
rect 66847 53065 66925 53111
rect 66971 53065 67049 53111
rect 67095 53065 67173 53111
rect 67219 53065 67297 53111
rect 67343 53065 67421 53111
rect 67467 53065 67545 53111
rect 67591 53065 67669 53111
rect 67715 53065 67793 53111
rect 67839 53065 67917 53111
rect 67963 53065 68041 53111
rect 68087 53065 68165 53111
rect 68211 53065 68289 53111
rect 68335 53065 68413 53111
rect 68459 53065 68537 53111
rect 68583 53065 68661 53111
rect 68707 53065 68785 53111
rect 68831 53065 68909 53111
rect 68955 53065 69033 53111
rect 69079 53065 69157 53111
rect 69203 53065 69281 53111
rect 69327 53065 69405 53111
rect 69451 53065 69529 53111
rect 69575 53065 69653 53111
rect 69699 53065 69777 53111
rect 69823 53065 69901 53111
rect 69947 53065 70025 53111
rect 70071 53065 70149 53111
rect 70195 53065 70273 53111
rect 70319 53065 70397 53111
rect 70443 53065 70521 53111
rect 70567 53065 70645 53111
rect 70691 53065 70769 53111
rect 70815 53065 70893 53111
rect 70939 53065 71017 53111
rect 71063 53065 71141 53111
rect 71187 53065 71265 53111
rect 71311 53065 71389 53111
rect 71435 53065 71513 53111
rect 71559 53065 71637 53111
rect 71683 53065 71761 53111
rect 71807 53065 71885 53111
rect 71931 53065 72009 53111
rect 72055 53065 72133 53111
rect 72179 53065 72257 53111
rect 72303 53065 72381 53111
rect 72427 53065 72505 53111
rect 72551 53065 72629 53111
rect 72675 53065 72753 53111
rect 72799 53065 72877 53111
rect 72923 53065 73001 53111
rect 73047 53065 73125 53111
rect 73171 53065 73249 53111
rect 73295 53065 73373 53111
rect 73419 53065 73497 53111
rect 73543 53065 73621 53111
rect 73667 53065 73745 53111
rect 73791 53065 73869 53111
rect 73915 53065 73993 53111
rect 74039 53065 74117 53111
rect 74163 53065 74241 53111
rect 74287 53065 74365 53111
rect 74411 53065 74489 53111
rect 74535 53065 74613 53111
rect 74659 53065 74737 53111
rect 74783 53065 74861 53111
rect 74907 53065 74985 53111
rect 75031 53065 75109 53111
rect 75155 53065 75233 53111
rect 75279 53065 75357 53111
rect 75403 53065 75481 53111
rect 75527 53065 75605 53111
rect 75651 53065 75729 53111
rect 75775 53065 75853 53111
rect 75899 53065 75977 53111
rect 76023 53065 76101 53111
rect 76147 53065 76225 53111
rect 76271 53065 76349 53111
rect 76395 53065 76473 53111
rect 76519 53065 76597 53111
rect 76643 53065 76721 53111
rect 76767 53065 76845 53111
rect 76891 53065 76969 53111
rect 77015 53065 77093 53111
rect 77139 53065 77217 53111
rect 77263 53065 77341 53111
rect 77387 53065 77465 53111
rect 77511 53065 77589 53111
rect 77635 53065 77713 53111
rect 77759 53065 77837 53111
rect 77883 53065 77961 53111
rect 78007 53065 78085 53111
rect 78131 53065 78209 53111
rect 78255 53065 78333 53111
rect 78379 53065 78457 53111
rect 78503 53065 78581 53111
rect 78627 53065 78705 53111
rect 78751 53065 78829 53111
rect 78875 53065 78953 53111
rect 78999 53065 79077 53111
rect 79123 53065 79201 53111
rect 79247 53065 79325 53111
rect 79371 53065 79449 53111
rect 79495 53065 79573 53111
rect 79619 53065 79697 53111
rect 79743 53065 79821 53111
rect 79867 53065 79945 53111
rect 79991 53065 80069 53111
rect 80115 53065 80193 53111
rect 80239 53065 80317 53111
rect 80363 53065 80441 53111
rect 80487 53065 80565 53111
rect 80611 53065 80689 53111
rect 80735 53065 80813 53111
rect 80859 53065 80937 53111
rect 80983 53065 81061 53111
rect 81107 53065 81185 53111
rect 81231 53065 81309 53111
rect 81355 53065 81433 53111
rect 81479 53065 81557 53111
rect 81603 53065 81681 53111
rect 81727 53065 81805 53111
rect 81851 53065 81929 53111
rect 81975 53065 82053 53111
rect 82099 53065 82177 53111
rect 82223 53065 82301 53111
rect 82347 53065 82425 53111
rect 82471 53065 82549 53111
rect 82595 53065 82673 53111
rect 82719 53065 82797 53111
rect 82843 53065 82921 53111
rect 82967 53065 83045 53111
rect 83091 53065 83169 53111
rect 83215 53065 83293 53111
rect 83339 53065 83417 53111
rect 83463 53065 83541 53111
rect 83587 53065 83665 53111
rect 83711 53065 83789 53111
rect 83835 53065 83913 53111
rect 83959 53065 84037 53111
rect 84083 53065 84161 53111
rect 84207 53065 84285 53111
rect 84331 53065 84409 53111
rect 84455 53065 84533 53111
rect 84579 53065 84657 53111
rect 84703 53065 84781 53111
rect 84827 53065 84905 53111
rect 84951 53065 85029 53111
rect 85075 53065 85153 53111
rect 85199 53065 85277 53111
rect 85323 53065 85401 53111
rect 85447 53065 85525 53111
rect 85571 53065 85649 53111
rect 85695 53065 85706 53111
rect 0 53054 85706 53065
rect 0 52963 1000 53054
rect 0 1117 89 52963
rect 435 1117 1000 52963
rect 0 1026 1000 1117
rect 85440 52963 85808 52974
rect 85440 1117 85451 52963
rect 85797 1117 85808 52963
rect 85440 1106 85808 1117
rect 0 1015 85706 1026
rect 0 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85706 1015
rect 0 891 85706 969
rect 0 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85706 891
rect 0 767 85706 845
rect 0 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85706 767
rect 0 643 85706 721
rect 0 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85706 643
rect 0 586 85706 597
rect 0 403 1000 586
<< metal2 >>
rect 424 403 1424 52949
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105905487112_128x8m81  M1_PSUB43105905487112_128x8m81_0
timestamp 1750858719
transform -1 0 85672 0 1 53088
box 0 0 1 1
use M1_PSUB43105905487112_128x8m81  M1_PSUB43105905487112_128x8m81_1
timestamp 1750858719
transform -1 0 85672 0 1 620
box 0 0 1 1
use M1_PSUB43105905487113_128x8m81  M1_PSUB43105905487113_128x8m81_0
timestamp 1750858719
transform 1 0 85474 0 1 1140
box 0 0 1 1
use M1_PSUB43105905487113_128x8m81  M1_PSUB43105905487113_128x8m81_1
timestamp 1750858719
transform 1 0 112 0 1 1140
box 0 0 1 1
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2235432
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2234776
string path 4.620 11.160 4.620 0.000 
<< end >>
