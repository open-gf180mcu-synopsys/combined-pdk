magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 5350 1094
<< pwell >>
rect -86 -86 5350 453
<< mvnmos >>
rect 124 69 244 333
rect 308 69 428 333
rect 532 69 652 333
rect 716 69 836 333
rect 940 69 1060 333
rect 1124 69 1244 333
rect 1348 69 1468 333
rect 1532 69 1652 333
rect 1890 69 2010 333
rect 2084 69 2204 333
rect 2308 69 2428 333
rect 2492 69 2612 333
rect 2716 69 2836 333
rect 2900 69 3020 333
rect 3124 69 3244 333
rect 3308 69 3428 333
rect 3532 69 3652 333
rect 3716 69 3836 333
rect 3940 69 4060 333
rect 4124 69 4244 333
rect 4348 69 4468 333
rect 4532 69 4652 333
rect 4756 69 4876 333
rect 4940 69 5060 333
<< mvpmos >>
rect 124 573 224 939
rect 328 573 428 939
rect 532 573 632 939
rect 736 573 836 939
rect 940 573 1040 939
rect 1144 573 1244 939
rect 1348 573 1448 939
rect 1552 573 1652 939
rect 1900 573 2000 939
rect 2104 573 2204 939
rect 2308 573 2408 939
rect 2512 573 2612 939
rect 2716 573 2816 939
rect 2920 573 3020 939
rect 3124 573 3224 939
rect 3328 573 3428 939
rect 3532 573 3632 939
rect 3736 573 3836 939
rect 3940 573 4040 939
rect 4144 573 4244 939
rect 4348 573 4448 939
rect 4552 573 4652 939
rect 4756 573 4856 939
rect 4960 573 5060 939
<< mvndiff >>
rect 36 239 124 333
rect 36 193 49 239
rect 95 193 124 239
rect 36 69 124 193
rect 244 69 308 333
rect 428 136 532 333
rect 428 90 457 136
rect 503 90 532 136
rect 428 69 532 90
rect 652 69 716 333
rect 836 239 940 333
rect 836 193 865 239
rect 911 193 940 239
rect 836 69 940 193
rect 1060 69 1124 333
rect 1244 136 1348 333
rect 1244 90 1273 136
rect 1319 90 1348 136
rect 1244 69 1348 90
rect 1468 69 1532 333
rect 1652 239 1890 333
rect 1652 193 1681 239
rect 1727 193 1890 239
rect 1652 69 1890 193
rect 2010 69 2084 333
rect 2204 136 2308 333
rect 2204 90 2233 136
rect 2279 90 2308 136
rect 2204 69 2308 90
rect 2428 69 2492 333
rect 2612 228 2716 333
rect 2612 182 2641 228
rect 2687 182 2716 228
rect 2612 69 2716 182
rect 2836 69 2900 333
rect 3020 128 3124 333
rect 3020 82 3049 128
rect 3095 82 3124 128
rect 3020 69 3124 82
rect 3244 69 3308 333
rect 3428 242 3532 333
rect 3428 196 3457 242
rect 3503 196 3532 242
rect 3428 69 3532 196
rect 3652 69 3716 333
rect 3836 128 3940 333
rect 3836 82 3865 128
rect 3911 82 3940 128
rect 3836 69 3940 82
rect 4060 69 4124 333
rect 4244 239 4348 333
rect 4244 193 4273 239
rect 4319 193 4348 239
rect 4244 69 4348 193
rect 4468 69 4532 333
rect 4652 128 4756 333
rect 4652 82 4681 128
rect 4727 82 4756 128
rect 4652 69 4756 82
rect 4876 69 4940 333
rect 5060 239 5148 333
rect 5060 193 5089 239
rect 5135 193 5148 239
rect 5060 69 5148 193
<< mvpdiff >>
rect 36 800 124 939
rect 36 660 49 800
rect 95 660 124 800
rect 36 573 124 660
rect 224 800 328 939
rect 224 660 253 800
rect 299 660 328 800
rect 224 573 328 660
rect 428 892 532 939
rect 428 752 457 892
rect 503 752 532 892
rect 428 573 532 752
rect 632 800 736 939
rect 632 660 661 800
rect 707 660 736 800
rect 632 573 736 660
rect 836 892 940 939
rect 836 752 865 892
rect 911 752 940 892
rect 836 573 940 752
rect 1040 800 1144 939
rect 1040 660 1069 800
rect 1115 660 1144 800
rect 1040 573 1144 660
rect 1244 863 1348 939
rect 1244 723 1273 863
rect 1319 723 1348 863
rect 1244 573 1348 723
rect 1448 800 1552 939
rect 1448 660 1477 800
rect 1523 660 1552 800
rect 1448 573 1552 660
rect 1652 860 1740 939
rect 1652 720 1681 860
rect 1727 720 1740 860
rect 1652 573 1740 720
rect 1812 860 1900 939
rect 1812 720 1825 860
rect 1871 720 1900 860
rect 1812 573 1900 720
rect 2000 769 2104 939
rect 2000 629 2029 769
rect 2075 629 2104 769
rect 2000 573 2104 629
rect 2204 861 2308 939
rect 2204 721 2233 861
rect 2279 721 2308 861
rect 2204 573 2308 721
rect 2408 769 2512 939
rect 2408 629 2437 769
rect 2483 629 2512 769
rect 2408 573 2512 629
rect 2612 861 2716 939
rect 2612 721 2641 861
rect 2687 721 2716 861
rect 2612 573 2716 721
rect 2816 769 2920 939
rect 2816 629 2845 769
rect 2891 629 2920 769
rect 2816 573 2920 629
rect 3020 843 3124 939
rect 3020 703 3049 843
rect 3095 703 3124 843
rect 3020 573 3124 703
rect 3224 769 3328 939
rect 3224 629 3253 769
rect 3299 629 3328 769
rect 3224 573 3328 629
rect 3428 832 3532 939
rect 3428 692 3457 832
rect 3503 692 3532 832
rect 3428 573 3532 692
rect 3632 769 3736 939
rect 3632 629 3661 769
rect 3707 629 3736 769
rect 3632 573 3736 629
rect 3836 843 3940 939
rect 3836 703 3865 843
rect 3911 703 3940 843
rect 3836 573 3940 703
rect 4040 769 4144 939
rect 4040 629 4069 769
rect 4115 629 4144 769
rect 4040 573 4144 629
rect 4244 861 4348 939
rect 4244 721 4273 861
rect 4319 721 4348 861
rect 4244 573 4348 721
rect 4448 769 4552 939
rect 4448 629 4477 769
rect 4523 629 4552 769
rect 4448 573 4552 629
rect 4652 843 4756 939
rect 4652 703 4681 843
rect 4727 703 4756 843
rect 4652 573 4756 703
rect 4856 769 4960 939
rect 4856 629 4885 769
rect 4931 629 4960 769
rect 4856 573 4960 629
rect 5060 800 5148 939
rect 5060 660 5089 800
rect 5135 660 5148 800
rect 5060 573 5148 660
<< mvndiffc >>
rect 49 193 95 239
rect 457 90 503 136
rect 865 193 911 239
rect 1273 90 1319 136
rect 1681 193 1727 239
rect 2233 90 2279 136
rect 2641 182 2687 228
rect 3049 82 3095 128
rect 3457 196 3503 242
rect 3865 82 3911 128
rect 4273 193 4319 239
rect 4681 82 4727 128
rect 5089 193 5135 239
<< mvpdiffc >>
rect 49 660 95 800
rect 253 660 299 800
rect 457 752 503 892
rect 661 660 707 800
rect 865 752 911 892
rect 1069 660 1115 800
rect 1273 723 1319 863
rect 1477 660 1523 800
rect 1681 720 1727 860
rect 1825 720 1871 860
rect 2029 629 2075 769
rect 2233 721 2279 861
rect 2437 629 2483 769
rect 2641 721 2687 861
rect 2845 629 2891 769
rect 3049 703 3095 843
rect 3253 629 3299 769
rect 3457 692 3503 832
rect 3661 629 3707 769
rect 3865 703 3911 843
rect 4069 629 4115 769
rect 4273 721 4319 861
rect 4477 629 4523 769
rect 4681 703 4727 843
rect 4885 629 4931 769
rect 5089 660 5135 800
<< polysilicon >>
rect 124 939 224 983
rect 328 939 428 983
rect 532 939 632 983
rect 736 939 836 983
rect 940 939 1040 983
rect 1144 939 1244 983
rect 1348 939 1448 983
rect 1552 939 1652 983
rect 1900 939 2000 983
rect 2104 939 2204 983
rect 2308 939 2408 983
rect 2512 939 2612 983
rect 2716 939 2816 983
rect 2920 939 3020 983
rect 3124 939 3224 983
rect 3328 939 3428 983
rect 3532 939 3632 983
rect 3736 939 3836 983
rect 3940 939 4040 983
rect 4144 939 4244 983
rect 4348 939 4448 983
rect 4552 939 4652 983
rect 4756 939 4856 983
rect 4960 939 5060 983
rect 124 500 224 573
rect 124 454 165 500
rect 211 454 224 500
rect 124 377 224 454
rect 328 513 428 573
rect 532 513 632 573
rect 328 500 632 513
rect 328 454 366 500
rect 412 454 632 500
rect 328 441 632 454
rect 328 377 428 441
rect 124 333 244 377
rect 308 333 428 377
rect 532 377 632 441
rect 736 513 836 573
rect 940 513 1040 573
rect 736 500 1040 513
rect 736 454 749 500
rect 795 454 1040 500
rect 736 441 1040 454
rect 736 377 836 441
rect 532 333 652 377
rect 716 333 836 377
rect 940 377 1040 441
rect 1144 513 1244 573
rect 1348 513 1448 573
rect 1144 500 1448 513
rect 1144 454 1157 500
rect 1203 454 1448 500
rect 1144 441 1448 454
rect 1144 377 1244 441
rect 940 333 1060 377
rect 1124 333 1244 377
rect 1348 377 1448 441
rect 1552 500 1652 573
rect 1552 454 1565 500
rect 1611 454 1652 500
rect 1552 377 1652 454
rect 1900 500 2000 573
rect 1900 454 1940 500
rect 1986 454 2000 500
rect 1900 377 2000 454
rect 2104 513 2204 573
rect 2308 513 2408 573
rect 2104 500 2408 513
rect 2104 454 2349 500
rect 2395 454 2408 500
rect 2104 441 2408 454
rect 2104 377 2204 441
rect 1348 333 1468 377
rect 1532 333 1652 377
rect 1890 333 2010 377
rect 2084 333 2204 377
rect 2308 377 2408 441
rect 2512 513 2612 573
rect 2716 513 2816 573
rect 2512 469 2816 513
rect 2512 423 2525 469
rect 2571 441 2816 469
rect 2571 423 2612 441
rect 2512 377 2612 423
rect 2308 333 2428 377
rect 2492 333 2612 377
rect 2716 377 2816 441
rect 2920 513 3020 573
rect 3124 513 3224 573
rect 3328 513 3428 573
rect 2920 500 3224 513
rect 2920 454 2933 500
rect 2979 454 3224 500
rect 2920 441 3224 454
rect 2920 377 3020 441
rect 2716 333 2836 377
rect 2900 333 3020 377
rect 3124 377 3224 441
rect 3308 500 3428 513
rect 3308 454 3321 500
rect 3367 454 3428 500
rect 3124 333 3244 377
rect 3308 333 3428 454
rect 3532 500 3632 573
rect 3532 454 3573 500
rect 3619 454 3632 500
rect 3532 377 3632 454
rect 3736 513 3836 573
rect 3940 513 4040 573
rect 3736 500 4040 513
rect 3736 454 3961 500
rect 4007 454 4040 500
rect 3736 441 4040 454
rect 3736 377 3836 441
rect 3532 333 3652 377
rect 3716 333 3836 377
rect 3940 377 4040 441
rect 4144 513 4244 573
rect 4348 513 4448 573
rect 4144 469 4448 513
rect 4144 423 4157 469
rect 4203 441 4448 469
rect 4203 423 4244 441
rect 4144 377 4244 423
rect 3940 333 4060 377
rect 4124 333 4244 377
rect 4348 377 4448 441
rect 4552 513 4652 573
rect 4756 513 4856 573
rect 4552 500 4856 513
rect 4552 454 4565 500
rect 4611 454 4856 500
rect 4552 441 4856 454
rect 4552 377 4652 441
rect 4348 333 4468 377
rect 4532 333 4652 377
rect 4756 377 4856 441
rect 4960 500 5060 573
rect 4960 454 4973 500
rect 5019 454 5060 500
rect 4960 377 5060 454
rect 4756 333 4876 377
rect 4940 333 5060 377
rect 124 25 244 69
rect 308 25 428 69
rect 532 25 652 69
rect 716 25 836 69
rect 940 25 1060 69
rect 1124 25 1244 69
rect 1348 25 1468 69
rect 1532 25 1652 69
rect 1890 25 2010 69
rect 2084 25 2204 69
rect 2308 25 2428 69
rect 2492 25 2612 69
rect 2716 25 2836 69
rect 2900 25 3020 69
rect 3124 25 3244 69
rect 3308 25 3428 69
rect 3532 25 3652 69
rect 3716 25 3836 69
rect 3940 25 4060 69
rect 4124 25 4244 69
rect 4348 25 4468 69
rect 4532 25 4652 69
rect 4756 25 4876 69
rect 4940 25 5060 69
<< polycontact >>
rect 165 454 211 500
rect 366 454 412 500
rect 749 454 795 500
rect 1157 454 1203 500
rect 1565 454 1611 500
rect 1940 454 1986 500
rect 2349 454 2395 500
rect 2525 423 2571 469
rect 2933 454 2979 500
rect 3321 454 3367 500
rect 3573 454 3619 500
rect 3961 454 4007 500
rect 4157 423 4203 469
rect 4565 454 4611 500
rect 4973 454 5019 500
<< metal1 >>
rect 0 918 5264 1098
rect 49 800 95 918
rect 457 892 503 918
rect 49 649 95 660
rect 253 800 299 811
rect 865 892 911 918
rect 457 741 503 752
rect 661 800 707 811
rect 299 660 661 695
rect 1273 863 1319 918
rect 865 741 911 752
rect 1069 800 1115 811
rect 707 660 1069 695
rect 1681 860 1727 918
rect 1273 712 1319 723
rect 1477 800 1523 811
rect 1115 663 1230 695
rect 1115 660 1477 663
rect 1681 709 1727 720
rect 1825 861 5135 872
rect 1825 860 2233 861
rect 1871 826 2233 860
rect 1825 709 1871 720
rect 2029 769 2075 780
rect 1881 663 2029 664
rect 1523 660 2029 663
rect 253 649 2029 660
rect 1186 629 2029 649
rect 2279 826 2641 861
rect 2233 710 2279 721
rect 2437 769 2483 780
rect 2075 629 2437 664
rect 2687 843 4273 861
rect 2687 826 3049 843
rect 2641 710 2687 721
rect 2845 769 2902 780
rect 2483 629 2845 664
rect 2891 646 2902 769
rect 3095 832 3865 843
rect 3095 826 3457 832
rect 3049 692 3095 703
rect 3253 769 3299 780
rect 2891 629 3253 646
rect 3503 826 3865 832
rect 3457 681 3503 692
rect 3661 769 3707 780
rect 1186 618 3299 629
rect 1186 617 1891 618
rect 657 571 1142 603
rect 2865 600 3299 618
rect 3533 629 3661 646
rect 3911 826 4273 843
rect 3865 692 3911 703
rect 4069 769 4115 780
rect 3948 646 4069 664
rect 3707 629 4069 646
rect 4319 843 5135 861
rect 4319 826 4681 843
rect 4273 710 4319 721
rect 4477 769 4523 780
rect 4115 629 4477 664
rect 4727 826 5135 843
rect 5089 800 5135 826
rect 4681 692 4727 703
rect 4885 769 4931 780
rect 4523 646 4644 664
rect 4523 629 4885 646
rect 5089 649 5135 660
rect 3533 618 4931 629
rect 3533 603 3985 618
rect 3457 600 3985 603
rect 4607 600 4931 618
rect 657 557 1203 571
rect 165 500 211 511
rect 165 397 211 454
rect 366 500 418 542
rect 412 489 418 500
rect 657 489 703 557
rect 1098 525 1203 557
rect 412 454 703 489
rect 366 443 703 454
rect 749 500 795 511
rect 749 397 795 454
rect 1157 500 1203 525
rect 2420 554 2828 572
rect 3457 557 3579 600
rect 2420 526 2979 554
rect 1157 443 1203 454
rect 1565 500 1611 511
rect 1565 430 1611 454
rect 1262 397 1611 430
rect 165 351 1611 397
rect 1934 500 1986 511
rect 2420 500 2466 526
rect 2791 508 2979 526
rect 1934 454 1940 500
rect 1934 320 1986 454
rect 2338 454 2349 500
rect 2395 454 2466 500
rect 2933 500 2979 508
rect 2338 366 2466 454
rect 2525 469 2571 480
rect 2933 443 2979 454
rect 3321 500 3367 511
rect 2525 331 2571 423
rect 3321 331 3367 454
rect 2525 320 3367 331
rect 1934 285 3367 320
rect 1934 274 2555 285
rect 3457 242 3503 557
rect 4027 554 4556 572
rect 3950 526 4611 554
rect 3573 500 3619 511
rect 3950 500 4064 526
rect 3950 454 3961 500
rect 4007 454 4064 500
rect 4519 500 4611 526
rect 4157 469 4203 480
rect 3573 430 3619 454
rect 3573 397 3890 430
rect 4519 454 4565 500
rect 4519 443 4611 454
rect 4973 500 5019 511
rect 4157 397 4203 423
rect 4973 397 5019 454
rect 3573 351 5019 397
rect 38 193 49 239
rect 95 193 865 239
rect 911 193 1681 239
rect 1727 228 1738 239
rect 2681 228 3457 231
rect 1727 193 2641 228
rect 38 182 2641 193
rect 2687 196 3457 228
rect 3503 196 4273 239
rect 2687 193 4273 196
rect 4319 193 5089 239
rect 5135 193 5146 239
rect 2687 185 5146 193
rect 2687 182 2698 185
rect 4946 142 5146 185
rect 446 90 457 136
rect 503 90 514 136
rect 1262 90 1273 136
rect 1319 90 1330 136
rect 2222 90 2233 136
rect 2279 90 2290 136
rect 3049 128 3095 139
rect 0 82 3049 90
rect 3865 128 3911 139
rect 3095 82 3865 90
rect 4681 128 4727 139
rect 3911 82 4681 90
rect 4727 82 5264 90
rect 0 -90 5264 82
<< labels >>
flabel metal1 s 4973 480 5019 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 4027 554 4556 572 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 3321 480 3367 511 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 2420 554 2828 572 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 1565 430 1611 511 0 FreeSans 200 0 0 0 C1
port 5 nsew default input
flabel metal1 s 657 571 1142 603 0 FreeSans 200 0 0 0 C2
port 6 nsew default input
flabel metal1 s 0 918 5264 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 4681 136 4727 139 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 4885 664 4931 780 0 FreeSans 200 0 0 0 ZN
port 7 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 3573 480 3619 511 1 A1
port 1 nsew default input
rlabel metal1 s 4973 430 5019 480 1 A1
port 1 nsew default input
rlabel metal1 s 4157 430 4203 480 1 A1
port 1 nsew default input
rlabel metal1 s 3573 430 3619 480 1 A1
port 1 nsew default input
rlabel metal1 s 4973 397 5019 430 1 A1
port 1 nsew default input
rlabel metal1 s 4157 397 4203 430 1 A1
port 1 nsew default input
rlabel metal1 s 3573 397 3890 430 1 A1
port 1 nsew default input
rlabel metal1 s 3573 351 5019 397 1 A1
port 1 nsew default input
rlabel metal1 s 3950 526 4611 554 1 A2
port 2 nsew default input
rlabel metal1 s 4519 454 4611 526 1 A2
port 2 nsew default input
rlabel metal1 s 3950 454 4064 526 1 A2
port 2 nsew default input
rlabel metal1 s 4519 443 4611 454 1 A2
port 2 nsew default input
rlabel metal1 s 1934 480 1986 511 1 B1
port 3 nsew default input
rlabel metal1 s 3321 331 3367 480 1 B1
port 3 nsew default input
rlabel metal1 s 2525 331 2571 480 1 B1
port 3 nsew default input
rlabel metal1 s 1934 331 1986 480 1 B1
port 3 nsew default input
rlabel metal1 s 2525 320 3367 331 1 B1
port 3 nsew default input
rlabel metal1 s 1934 320 1986 331 1 B1
port 3 nsew default input
rlabel metal1 s 1934 285 3367 320 1 B1
port 3 nsew default input
rlabel metal1 s 1934 274 2555 285 1 B1
port 3 nsew default input
rlabel metal1 s 2420 526 2979 554 1 B2
port 4 nsew default input
rlabel metal1 s 2791 508 2979 526 1 B2
port 4 nsew default input
rlabel metal1 s 2420 508 2466 526 1 B2
port 4 nsew default input
rlabel metal1 s 2933 500 2979 508 1 B2
port 4 nsew default input
rlabel metal1 s 2420 500 2466 508 1 B2
port 4 nsew default input
rlabel metal1 s 2933 443 2979 500 1 B2
port 4 nsew default input
rlabel metal1 s 2338 443 2466 500 1 B2
port 4 nsew default input
rlabel metal1 s 2338 366 2466 443 1 B2
port 4 nsew default input
rlabel metal1 s 749 430 795 511 1 C1
port 5 nsew default input
rlabel metal1 s 165 430 211 511 1 C1
port 5 nsew default input
rlabel metal1 s 1262 397 1611 430 1 C1
port 5 nsew default input
rlabel metal1 s 749 397 795 430 1 C1
port 5 nsew default input
rlabel metal1 s 165 397 211 430 1 C1
port 5 nsew default input
rlabel metal1 s 165 351 1611 397 1 C1
port 5 nsew default input
rlabel metal1 s 657 557 1203 571 1 C2
port 6 nsew default input
rlabel metal1 s 1098 542 1203 557 1 C2
port 6 nsew default input
rlabel metal1 s 657 542 703 557 1 C2
port 6 nsew default input
rlabel metal1 s 1098 525 1203 542 1 C2
port 6 nsew default input
rlabel metal1 s 657 525 703 542 1 C2
port 6 nsew default input
rlabel metal1 s 366 525 418 542 1 C2
port 6 nsew default input
rlabel metal1 s 1157 489 1203 525 1 C2
port 6 nsew default input
rlabel metal1 s 657 489 703 525 1 C2
port 6 nsew default input
rlabel metal1 s 366 489 418 525 1 C2
port 6 nsew default input
rlabel metal1 s 1157 443 1203 489 1 C2
port 6 nsew default input
rlabel metal1 s 366 443 703 489 1 C2
port 6 nsew default input
rlabel metal1 s 4477 664 4523 780 1 ZN
port 7 nsew default output
rlabel metal1 s 4069 664 4115 780 1 ZN
port 7 nsew default output
rlabel metal1 s 3661 664 3707 780 1 ZN
port 7 nsew default output
rlabel metal1 s 4885 646 4931 664 1 ZN
port 7 nsew default output
rlabel metal1 s 3948 646 4644 664 1 ZN
port 7 nsew default output
rlabel metal1 s 3661 646 3707 664 1 ZN
port 7 nsew default output
rlabel metal1 s 3533 618 4931 646 1 ZN
port 7 nsew default output
rlabel metal1 s 4607 603 4931 618 1 ZN
port 7 nsew default output
rlabel metal1 s 3533 603 3985 618 1 ZN
port 7 nsew default output
rlabel metal1 s 4607 600 4931 603 1 ZN
port 7 nsew default output
rlabel metal1 s 3457 600 3985 603 1 ZN
port 7 nsew default output
rlabel metal1 s 3457 557 3579 600 1 ZN
port 7 nsew default output
rlabel metal1 s 3457 239 3503 557 1 ZN
port 7 nsew default output
rlabel metal1 s 3457 231 5146 239 1 ZN
port 7 nsew default output
rlabel metal1 s 38 231 1738 239 1 ZN
port 7 nsew default output
rlabel metal1 s 2681 228 5146 231 1 ZN
port 7 nsew default output
rlabel metal1 s 38 228 1738 231 1 ZN
port 7 nsew default output
rlabel metal1 s 38 185 5146 228 1 ZN
port 7 nsew default output
rlabel metal1 s 4946 182 5146 185 1 ZN
port 7 nsew default output
rlabel metal1 s 38 182 2698 185 1 ZN
port 7 nsew default output
rlabel metal1 s 4946 142 5146 182 1 ZN
port 7 nsew default output
rlabel metal1 s 1681 741 1727 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1273 741 1319 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 865 741 911 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 457 741 503 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 741 95 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1681 712 1727 741 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1273 712 1319 741 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 712 95 741 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1681 709 1727 712 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 709 95 712 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 649 95 709 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3865 136 3911 139 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3049 136 3095 139 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 4681 90 4727 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3865 90 3911 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3049 90 3095 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 2222 90 2290 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1262 90 1330 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 446 90 514 136 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5264 90 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5264 1008
string GDS_END 1258708
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1247576
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
