magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1720 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 850 210 910 380
rect 1020 210 1080 380
rect 1240 210 1300 380
rect 1410 210 1470 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
rect 850 720 910 1060
rect 1020 720 1080 1060
rect 1240 720 1300 1060
rect 1410 720 1470 1060
<< ndiff >>
rect 90 298 190 380
rect 90 252 112 298
rect 158 252 190 298
rect 90 210 190 252
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 530 380
rect 590 318 690 380
rect 590 272 622 318
rect 668 272 690 318
rect 590 210 690 272
rect 750 283 850 380
rect 750 237 772 283
rect 818 237 850 283
rect 750 210 850 237
rect 910 358 1020 380
rect 910 312 942 358
rect 988 312 1020 358
rect 910 210 1020 312
rect 1080 283 1240 380
rect 1080 237 1112 283
rect 1158 237 1240 283
rect 1080 210 1240 237
rect 1300 318 1410 380
rect 1300 272 1332 318
rect 1378 272 1410 318
rect 1300 210 1410 272
rect 1470 318 1620 380
rect 1470 272 1552 318
rect 1598 272 1620 318
rect 1470 210 1620 272
<< pdiff >>
rect 90 1032 190 1060
rect 90 798 112 1032
rect 158 798 190 1032
rect 90 720 190 798
rect 250 1007 360 1060
rect 250 773 282 1007
rect 328 773 360 1007
rect 250 720 360 773
rect 420 1007 530 1060
rect 420 773 452 1007
rect 498 773 530 1007
rect 420 720 530 773
rect 590 1007 690 1060
rect 590 773 622 1007
rect 668 773 690 1007
rect 590 720 690 773
rect 750 1007 850 1060
rect 750 773 772 1007
rect 818 773 850 1007
rect 750 720 850 773
rect 910 720 1020 1060
rect 1080 1007 1240 1060
rect 1080 773 1137 1007
rect 1183 773 1240 1007
rect 1080 720 1240 773
rect 1300 1013 1410 1060
rect 1300 967 1332 1013
rect 1378 967 1410 1013
rect 1300 720 1410 967
rect 1470 1007 1620 1060
rect 1470 773 1527 1007
rect 1573 773 1620 1007
rect 1470 720 1620 773
<< ndiffc >>
rect 112 252 158 298
rect 282 272 328 318
rect 622 272 668 318
rect 772 237 818 283
rect 942 312 988 358
rect 1112 237 1158 283
rect 1332 272 1378 318
rect 1552 272 1598 318
<< pdiffc >>
rect 112 798 158 1032
rect 282 773 328 1007
rect 452 773 498 1007
rect 622 773 668 1007
rect 772 773 818 1007
rect 1137 773 1183 1007
rect 1332 967 1378 1013
rect 1527 773 1573 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1310 118 1460 140
rect 1310 72 1362 118
rect 1408 72 1460 118
rect 1310 50 1460 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1362 72 1408 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 850 1060 910 1110
rect 1020 1060 1080 1110
rect 1240 1060 1300 1110
rect 1410 1060 1470 1110
rect 190 690 250 720
rect 190 663 310 690
rect 190 617 237 663
rect 283 617 310 663
rect 190 590 310 617
rect 190 380 250 590
rect 360 540 420 720
rect 300 513 420 540
rect 530 530 590 720
rect 850 540 910 720
rect 300 467 327 513
rect 373 467 420 513
rect 300 440 420 467
rect 360 380 420 440
rect 470 503 590 530
rect 470 457 497 503
rect 543 457 590 503
rect 470 430 590 457
rect 780 513 910 540
rect 780 467 807 513
rect 853 467 910 513
rect 780 440 910 467
rect 530 380 590 430
rect 850 380 910 440
rect 1020 500 1080 720
rect 1240 700 1300 720
rect 1240 673 1360 700
rect 1240 627 1287 673
rect 1333 627 1360 673
rect 1240 600 1360 627
rect 1020 473 1120 500
rect 1020 427 1047 473
rect 1093 427 1120 473
rect 1020 400 1120 427
rect 1020 380 1080 400
rect 1240 380 1300 600
rect 1410 540 1470 720
rect 1350 513 1470 540
rect 1350 467 1377 513
rect 1423 467 1470 513
rect 1350 440 1470 467
rect 1410 380 1470 440
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 850 160 910 210
rect 1020 160 1080 210
rect 1240 160 1300 210
rect 1410 160 1470 210
<< polycontact >>
rect 237 617 283 663
rect 327 467 373 513
rect 497 457 543 503
rect 807 467 853 513
rect 1287 627 1333 673
rect 1047 427 1093 473
rect 1377 467 1423 513
<< metal1 >>
rect 0 1198 1720 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1720 1198
rect 0 1130 1720 1152
rect 110 1032 160 1060
rect 110 798 112 1032
rect 158 798 160 1032
rect 110 780 160 798
rect 280 1007 330 1130
rect 80 776 180 780
rect 80 724 104 776
rect 156 724 180 776
rect 80 720 180 724
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 720 330 773
rect 450 1007 500 1060
rect 450 773 452 1007
rect 498 773 500 1007
rect 110 298 160 720
rect 450 670 500 773
rect 620 1007 670 1130
rect 620 773 622 1007
rect 668 773 670 1007
rect 620 720 670 773
rect 770 1007 820 1130
rect 770 773 772 1007
rect 818 773 820 1007
rect 770 720 820 773
rect 1110 1007 1210 1060
rect 1110 773 1137 1007
rect 1183 773 1210 1007
rect 1330 1013 1380 1130
rect 1330 967 1332 1013
rect 1378 967 1380 1013
rect 1330 920 1380 967
rect 1500 1007 1600 1060
rect 1110 720 1210 773
rect 1500 773 1527 1007
rect 1573 773 1600 1007
rect 1500 720 1600 773
rect 210 666 700 670
rect 210 663 624 666
rect 210 617 237 663
rect 283 617 624 663
rect 210 614 624 617
rect 676 614 700 666
rect 1110 620 1160 720
rect 1260 676 1360 680
rect 1260 624 1284 676
rect 1336 624 1360 676
rect 1550 660 1600 720
rect 1550 650 1620 660
rect 1260 620 1360 624
rect 1540 646 1640 650
rect 210 610 700 614
rect 300 516 400 520
rect 300 464 324 516
rect 376 464 400 516
rect 300 460 400 464
rect 470 503 570 510
rect 470 457 497 503
rect 543 457 570 503
rect 470 450 570 457
rect 490 390 550 450
rect 470 386 570 390
rect 110 252 112 298
rect 158 252 160 298
rect 110 210 160 252
rect 280 318 330 380
rect 470 334 494 386
rect 546 334 570 386
rect 470 330 570 334
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 620 318 670 610
rect 940 570 1210 620
rect 1540 594 1564 646
rect 1616 594 1640 646
rect 1540 590 1640 594
rect 1550 580 1620 590
rect 780 516 880 520
rect 780 464 804 516
rect 856 464 880 516
rect 780 460 880 464
rect 620 272 622 318
rect 668 272 670 318
rect 940 358 990 570
rect 1150 520 1350 570
rect 1300 513 1450 520
rect 1040 476 1100 500
rect 1040 424 1044 476
rect 1096 424 1100 476
rect 1300 467 1377 513
rect 1423 467 1450 513
rect 1300 460 1450 467
rect 1040 400 1100 424
rect 940 312 942 358
rect 988 312 990 358
rect 620 210 670 272
rect 770 283 820 310
rect 940 290 990 312
rect 1330 318 1380 380
rect 770 237 772 283
rect 818 240 820 283
rect 1110 283 1160 310
rect 1110 240 1112 283
rect 818 237 1112 240
rect 1158 237 1160 283
rect 770 190 1160 237
rect 1330 272 1332 318
rect 1378 272 1380 318
rect 1330 140 1380 272
rect 1550 318 1600 580
rect 1550 272 1552 318
rect 1598 272 1600 318
rect 1550 210 1600 272
rect 0 118 1720 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1362 118
rect 1408 72 1720 118
rect 0 0 1720 72
<< via1 >>
rect 104 724 156 776
rect 624 614 676 666
rect 1284 673 1336 676
rect 1284 627 1287 673
rect 1287 627 1333 673
rect 1333 627 1336 673
rect 1284 624 1336 627
rect 324 513 376 516
rect 324 467 327 513
rect 327 467 373 513
rect 373 467 376 513
rect 324 464 376 467
rect 494 334 546 386
rect 1564 594 1616 646
rect 804 513 856 516
rect 804 467 807 513
rect 807 467 853 513
rect 853 467 856 513
rect 804 464 856 467
rect 1044 473 1096 476
rect 1044 427 1047 473
rect 1047 427 1093 473
rect 1093 427 1096 473
rect 1044 424 1096 427
<< metal2 >>
rect 80 776 180 790
rect 80 724 104 776
rect 156 724 180 776
rect 80 710 180 724
rect 600 670 700 680
rect 1260 676 1360 690
rect 1260 670 1284 676
rect 600 666 1284 670
rect 600 614 624 666
rect 676 624 1284 666
rect 1336 624 1360 676
rect 676 614 1360 624
rect 600 610 1360 614
rect 1540 646 1640 660
rect 600 600 700 610
rect 1540 594 1564 646
rect 1616 594 1640 646
rect 1540 580 1640 594
rect 300 520 400 530
rect 780 520 880 530
rect 300 516 880 520
rect 300 464 324 516
rect 376 464 804 516
rect 856 464 880 516
rect 1040 490 1100 500
rect 300 460 880 464
rect 300 450 400 460
rect 780 450 880 460
rect 1030 476 1110 490
rect 1030 424 1044 476
rect 1096 424 1110 476
rect 1030 410 1110 424
rect 480 390 560 400
rect 1030 390 1100 410
rect 470 386 1100 390
rect 470 334 494 386
rect 546 334 1100 386
rect 470 330 1100 334
rect 480 320 560 330
<< labels >>
rlabel via1 s 804 464 856 516 4 A
port 1 nsew signal input
rlabel via1 s 1044 424 1096 476 4 B
port 2 nsew signal input
rlabel via1 s 1564 594 1616 646 4 S
port 3 nsew signal output
rlabel via1 s 104 724 156 776 4 CO
port 4 nsew signal output
rlabel metal1 s 280 720 330 1270 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 620 720 670 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 770 720 820 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1330 920 1380 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1720 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1330 0 1380 380 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1720 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel via1 s 324 464 376 516 1 A
port 1 nsew signal input
rlabel metal2 s 300 450 400 530 1 A
port 1 nsew signal input
rlabel metal2 s 300 460 880 520 1 A
port 1 nsew signal input
rlabel metal2 s 780 450 880 530 1 A
port 1 nsew signal input
rlabel metal1 s 300 460 400 520 1 A
port 1 nsew signal input
rlabel metal1 s 780 460 880 520 1 A
port 1 nsew signal input
rlabel via1 s 494 334 546 386 1 B
port 2 nsew signal input
rlabel metal2 s 480 320 560 400 1 B
port 2 nsew signal input
rlabel metal2 s 470 330 1100 390 1 B
port 2 nsew signal input
rlabel metal2 s 1030 330 1100 490 1 B
port 2 nsew signal input
rlabel metal2 s 1040 330 1100 500 1 B
port 2 nsew signal input
rlabel metal2 s 1030 410 1110 490 1 B
port 2 nsew signal input
rlabel metal1 s 490 330 550 510 1 B
port 2 nsew signal input
rlabel metal1 s 470 330 570 390 1 B
port 2 nsew signal input
rlabel metal1 s 470 450 570 510 1 B
port 2 nsew signal input
rlabel metal1 s 1040 400 1100 500 1 B
port 2 nsew signal input
rlabel metal2 s 80 710 180 790 1 CO
port 4 nsew signal output
rlabel metal1 s 110 210 160 1060 1 CO
port 4 nsew signal output
rlabel metal1 s 80 720 180 780 1 CO
port 4 nsew signal output
rlabel metal2 s 1540 580 1640 660 1 S
port 3 nsew signal output
rlabel metal1 s 1550 210 1600 1060 1 S
port 3 nsew signal output
rlabel metal1 s 1500 720 1600 1060 1 S
port 3 nsew signal output
rlabel metal1 s 1550 580 1620 660 1 S
port 3 nsew signal output
rlabel metal1 s 1540 590 1640 650 1 S
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1720 1270
string GDS_END 30928
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 19812
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
