magic
tech gf180mcuA
timestamp 1750858719
<< properties >>
string GDS_END 500660
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 498928
<< end >>
