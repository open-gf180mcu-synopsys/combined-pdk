//Verilog HDL for "ECE733", "inverter" "functional"


module gf180mcu_fd_sc_mcu7t5v0__inv_1 ( I, ZN, VDD, VSS );

  input I;
  output ZN;
  inout VDD;
  inout VSS;
  assign ZN = ~I;
endmodule
