magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 2900 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 570 210 630 380
rect 800 210 860 380
rect 910 210 970 380
rect 1080 210 1140 380
rect 1190 210 1250 380
rect 1420 210 1480 380
rect 1630 210 1690 380
rect 1800 210 1860 380
rect 2160 210 2220 380
rect 2480 210 2540 380
rect 2650 210 2710 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 570 720 630 1060
rect 800 720 860 1060
rect 910 720 970 1060
rect 1080 720 1140 1060
rect 1190 720 1250 1060
rect 1420 720 1480 1060
rect 1630 720 1690 1060
rect 1800 720 1860 1060
rect 2160 720 2220 1060
rect 2480 720 2540 1060
rect 2650 720 2710 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 283 360 380
rect 250 237 282 283
rect 328 237 360 283
rect 250 210 360 237
rect 420 210 570 380
rect 630 283 800 380
rect 630 237 692 283
rect 738 237 800 283
rect 630 210 800 237
rect 860 210 910 380
rect 970 278 1080 380
rect 970 232 1002 278
rect 1048 232 1080 278
rect 970 210 1080 232
rect 1140 210 1190 380
rect 1250 278 1420 380
rect 1250 232 1312 278
rect 1358 232 1420 278
rect 1250 210 1420 232
rect 1480 210 1630 380
rect 1690 283 1800 380
rect 1690 237 1722 283
rect 1768 237 1800 283
rect 1690 210 1800 237
rect 1860 278 1960 380
rect 1860 232 1892 278
rect 1938 232 1960 278
rect 1860 210 1960 232
rect 2060 278 2160 380
rect 2060 232 2082 278
rect 2128 232 2160 278
rect 2060 210 2160 232
rect 2220 318 2320 380
rect 2220 272 2252 318
rect 2298 272 2320 318
rect 2220 210 2320 272
rect 2380 318 2480 380
rect 2380 272 2402 318
rect 2448 272 2480 318
rect 2380 210 2480 272
rect 2540 298 2650 380
rect 2540 252 2572 298
rect 2618 252 2650 298
rect 2540 210 2650 252
rect 2710 318 2810 380
rect 2710 272 2742 318
rect 2788 272 2810 318
rect 2710 210 2810 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1038 360 1060
rect 250 992 282 1038
rect 328 992 360 1038
rect 250 720 360 992
rect 420 720 570 1060
rect 630 1030 800 1060
rect 630 890 692 1030
rect 738 890 800 1030
rect 630 720 800 890
rect 860 720 910 1060
rect 970 1020 1080 1060
rect 970 880 1002 1020
rect 1048 880 1080 1020
rect 970 720 1080 880
rect 1140 720 1190 1060
rect 1250 1030 1420 1060
rect 1250 890 1312 1030
rect 1358 890 1420 1030
rect 1250 720 1420 890
rect 1480 720 1630 1060
rect 1690 1038 1800 1060
rect 1690 992 1722 1038
rect 1768 992 1800 1038
rect 1690 720 1800 992
rect 1860 1007 1960 1060
rect 1860 773 1892 1007
rect 1938 773 1960 1007
rect 1860 720 1960 773
rect 2060 1007 2160 1060
rect 2060 773 2082 1007
rect 2128 773 2160 1007
rect 2060 720 2160 773
rect 2220 1007 2320 1060
rect 2220 773 2252 1007
rect 2298 773 2320 1007
rect 2220 720 2320 773
rect 2380 1007 2480 1060
rect 2380 773 2402 1007
rect 2448 773 2480 1007
rect 2380 720 2480 773
rect 2540 1015 2650 1060
rect 2540 875 2572 1015
rect 2618 875 2650 1015
rect 2540 720 2650 875
rect 2710 998 2810 1060
rect 2710 952 2742 998
rect 2788 952 2810 998
rect 2710 720 2810 952
<< ndiffc >>
rect 112 272 158 318
rect 282 237 328 283
rect 692 237 738 283
rect 1002 232 1048 278
rect 1312 232 1358 278
rect 1722 237 1768 283
rect 1892 232 1938 278
rect 2082 232 2128 278
rect 2252 272 2298 318
rect 2402 272 2448 318
rect 2572 252 2618 298
rect 2742 272 2788 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 992 328 1038
rect 692 890 738 1030
rect 1002 880 1048 1020
rect 1312 890 1358 1030
rect 1722 992 1768 1038
rect 1892 773 1938 1007
rect 2082 773 2128 1007
rect 2252 773 2298 1007
rect 2402 773 2448 1007
rect 2572 875 2618 1015
rect 2742 952 2788 998
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
rect 1500 1198 1650 1220
rect 1500 1152 1552 1198
rect 1598 1152 1650 1198
rect 1500 1130 1650 1152
rect 1740 1198 1890 1220
rect 1740 1152 1792 1198
rect 1838 1152 1890 1198
rect 1740 1130 1890 1152
rect 1980 1198 2130 1220
rect 1980 1152 2032 1198
rect 2078 1152 2130 1198
rect 1980 1130 2130 1152
rect 2220 1198 2370 1220
rect 2220 1152 2272 1198
rect 2318 1152 2370 1198
rect 2220 1130 2370 1152
rect 2460 1198 2610 1220
rect 2460 1152 2512 1198
rect 2558 1152 2610 1198
rect 2460 1130 2610 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
rect 1552 1152 1598 1198
rect 1792 1152 1838 1198
rect 2032 1152 2078 1198
rect 2272 1152 2318 1198
rect 2512 1152 2558 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 570 1060 630 1110
rect 800 1060 860 1110
rect 910 1060 970 1110
rect 1080 1060 1140 1110
rect 1190 1060 1250 1110
rect 1420 1060 1480 1110
rect 1630 1060 1690 1110
rect 1800 1060 1860 1110
rect 2160 1060 2220 1110
rect 2480 1060 2540 1110
rect 2650 1060 2710 1110
rect 190 700 250 720
rect 190 673 290 700
rect 190 627 217 673
rect 263 627 290 673
rect 360 670 420 720
rect 570 700 630 720
rect 500 678 630 700
rect 190 600 290 627
rect 340 643 450 670
rect 190 380 250 600
rect 340 597 377 643
rect 423 597 450 643
rect 500 632 532 678
rect 578 670 630 678
rect 578 632 600 670
rect 500 610 600 632
rect 340 570 450 597
rect 800 590 860 720
rect 910 700 970 720
rect 1080 700 1140 720
rect 910 630 1140 700
rect 360 380 420 570
rect 650 540 860 590
rect 650 500 710 540
rect 530 473 710 500
rect 990 490 1050 630
rect 1190 590 1250 720
rect 1420 700 1480 720
rect 1420 673 1540 700
rect 1420 670 1467 673
rect 1440 627 1467 670
rect 1513 627 1540 673
rect 1440 600 1540 627
rect 1190 540 1390 590
rect 1630 540 1690 720
rect 1800 670 1860 720
rect 1800 643 1900 670
rect 1800 597 1827 643
rect 1873 597 1900 643
rect 2160 610 2220 720
rect 2480 610 2540 720
rect 1800 570 1900 597
rect 2100 583 2220 610
rect 1340 520 1390 540
rect 530 427 567 473
rect 613 427 710 473
rect 530 420 710 427
rect 760 468 860 490
rect 760 422 787 468
rect 833 422 860 468
rect 530 400 650 420
rect 760 400 860 422
rect 570 380 630 400
rect 800 380 860 400
rect 910 480 1050 490
rect 910 468 1140 480
rect 910 422 947 468
rect 993 422 1140 468
rect 910 400 1140 422
rect 910 380 970 400
rect 1080 380 1140 400
rect 1190 468 1290 490
rect 1190 422 1217 468
rect 1263 422 1290 468
rect 1190 400 1290 422
rect 1340 473 1480 520
rect 1340 427 1397 473
rect 1443 427 1480 473
rect 1610 513 1710 540
rect 1610 467 1637 513
rect 1683 467 1710 513
rect 1610 440 1710 467
rect 1340 420 1480 427
rect 1370 400 1480 420
rect 1190 380 1250 400
rect 1420 380 1480 400
rect 1630 380 1690 440
rect 1800 380 1860 570
rect 2100 537 2127 583
rect 2173 537 2220 583
rect 2100 510 2220 537
rect 2430 583 2540 610
rect 2430 537 2457 583
rect 2503 537 2540 583
rect 2650 540 2710 720
rect 2430 510 2540 537
rect 2160 380 2220 510
rect 2480 380 2540 510
rect 2590 513 2710 540
rect 2590 467 2617 513
rect 2663 467 2710 513
rect 2590 440 2710 467
rect 2650 380 2710 440
rect 190 160 250 210
rect 360 160 420 210
rect 570 160 630 210
rect 800 160 860 210
rect 910 160 970 210
rect 1080 160 1140 210
rect 1190 160 1250 210
rect 1420 160 1480 210
rect 1630 160 1690 210
rect 1800 160 1860 210
rect 2160 160 2220 210
rect 2480 160 2540 210
rect 2650 160 2710 210
<< polycontact >>
rect 217 627 263 673
rect 377 597 423 643
rect 532 632 578 678
rect 1467 627 1513 673
rect 1827 597 1873 643
rect 567 427 613 473
rect 787 422 833 468
rect 947 422 993 468
rect 1217 422 1263 468
rect 1397 427 1443 473
rect 1637 467 1683 513
rect 2127 537 2173 583
rect 2457 537 2503 583
rect 2617 467 2663 513
<< metal1 >>
rect 0 1198 2900 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1552 1198
rect 1598 1152 1792 1198
rect 1838 1152 2032 1198
rect 2078 1152 2272 1198
rect 2318 1152 2512 1198
rect 2558 1152 2900 1198
rect 0 1130 2900 1152
rect 110 1007 160 1060
rect 110 773 112 1007
rect 158 773 160 1007
rect 280 1038 330 1130
rect 280 992 282 1038
rect 328 992 330 1038
rect 280 970 330 992
rect 660 1030 770 1060
rect 660 920 692 1030
rect 110 490 160 773
rect 100 480 160 490
rect 80 476 160 480
rect 80 424 104 476
rect 156 424 160 476
rect 80 420 160 424
rect 100 400 160 420
rect 110 318 160 400
rect 210 890 692 920
rect 738 890 770 1030
rect 210 860 770 890
rect 1000 1020 1050 1130
rect 1000 880 1002 1020
rect 1048 880 1050 1020
rect 210 680 270 860
rect 1000 840 1050 880
rect 1280 1030 1390 1060
rect 1280 916 1312 1030
rect 1280 864 1304 916
rect 1358 890 1390 1030
rect 1720 1038 1770 1130
rect 1720 992 1722 1038
rect 1768 992 1770 1038
rect 1720 970 1770 992
rect 1890 1007 1940 1060
rect 1356 864 1390 890
rect 1280 840 1390 864
rect 1610 916 1710 920
rect 1610 864 1634 916
rect 1686 864 1710 916
rect 1610 860 1710 864
rect 1630 840 1690 860
rect 1890 773 1892 1007
rect 1938 773 1940 1007
rect 1890 770 1940 773
rect 2080 1007 2130 1130
rect 2080 773 2082 1007
rect 2128 773 2130 1007
rect 1890 720 2000 770
rect 2080 720 2130 773
rect 2250 1007 2300 1060
rect 2250 773 2252 1007
rect 2298 773 2300 1007
rect 210 673 290 680
rect 210 627 217 673
rect 263 627 290 673
rect 500 678 1790 680
rect 210 620 290 627
rect 350 646 450 650
rect 210 430 270 620
rect 350 594 374 646
rect 426 594 450 646
rect 500 632 532 678
rect 578 673 1790 678
rect 578 632 1467 673
rect 500 627 1467 632
rect 1513 670 1790 673
rect 1513 650 1880 670
rect 1513 646 1900 650
rect 1513 627 1824 646
rect 500 620 1824 627
rect 350 590 450 594
rect 780 480 840 620
rect 940 480 1000 490
rect 540 476 640 480
rect 210 380 450 430
rect 540 424 564 476
rect 616 424 640 476
rect 540 420 640 424
rect 760 468 860 480
rect 760 422 787 468
rect 833 422 860 468
rect 760 420 860 422
rect 920 476 1020 480
rect 920 424 944 476
rect 996 424 1020 476
rect 1210 470 1270 620
rect 1800 594 1824 620
rect 1876 594 1900 646
rect 1800 590 1900 594
rect 1950 520 2000 720
rect 1610 516 1710 520
rect 1390 480 1450 500
rect 1380 473 1510 480
rect 920 422 947 424
rect 993 422 1020 424
rect 920 420 1020 422
rect 1190 468 1290 470
rect 1190 422 1217 468
rect 1263 422 1290 468
rect 1190 410 1290 422
rect 1380 427 1397 473
rect 1443 427 1510 473
rect 1610 464 1634 516
rect 1686 464 1710 516
rect 1610 460 1710 464
rect 1890 460 2000 520
rect 2120 583 2180 610
rect 2120 537 2127 583
rect 2173 537 2180 583
rect 1380 420 1510 427
rect 1390 400 1510 420
rect 400 350 450 380
rect 1450 386 1510 400
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 283 330 320
rect 400 300 770 350
rect 1280 346 1390 350
rect 280 237 282 283
rect 328 237 330 283
rect 280 140 330 237
rect 660 283 770 300
rect 660 237 692 283
rect 738 237 770 283
rect 660 210 770 237
rect 1000 278 1050 300
rect 1000 232 1002 278
rect 1048 232 1050 278
rect 1000 140 1050 232
rect 1280 294 1304 346
rect 1356 294 1390 346
rect 1450 334 1454 386
rect 1506 334 1510 386
rect 1450 310 1510 334
rect 1890 386 1950 460
rect 2120 410 2180 537
rect 2250 590 2300 773
rect 2400 1007 2450 1060
rect 2400 773 2402 1007
rect 2448 780 2450 1007
rect 2570 1015 2620 1130
rect 2570 875 2572 1015
rect 2618 875 2620 1015
rect 2570 830 2620 875
rect 2740 998 2790 1060
rect 2740 952 2742 998
rect 2788 952 2790 998
rect 2740 920 2790 952
rect 2740 906 2850 920
rect 2740 854 2774 906
rect 2826 854 2850 906
rect 2740 850 2850 854
rect 2740 840 2840 850
rect 2448 776 2690 780
rect 2448 773 2614 776
rect 2400 724 2614 773
rect 2666 724 2690 776
rect 2400 720 2690 724
rect 2250 586 2530 590
rect 2250 534 2454 586
rect 2506 534 2530 586
rect 2250 530 2530 534
rect 1890 334 1894 386
rect 1946 334 1950 386
rect 2100 406 2200 410
rect 2100 354 2124 406
rect 2176 354 2200 406
rect 2100 350 2200 354
rect 1280 278 1390 294
rect 1280 232 1312 278
rect 1358 232 1390 278
rect 1280 210 1390 232
rect 1720 283 1770 320
rect 1720 237 1722 283
rect 1768 237 1770 283
rect 1720 140 1770 237
rect 1890 310 1950 334
rect 2250 318 2300 530
rect 2610 513 2670 720
rect 2610 467 2617 513
rect 2663 467 2670 513
rect 2610 440 2670 467
rect 1890 278 1940 310
rect 1890 232 1892 278
rect 1938 232 1940 278
rect 1890 210 1940 232
rect 2080 278 2130 300
rect 2080 232 2082 278
rect 2128 232 2130 278
rect 2080 140 2130 232
rect 2250 272 2252 318
rect 2298 272 2300 318
rect 2250 210 2300 272
rect 2400 390 2670 440
rect 2400 318 2450 390
rect 2400 272 2402 318
rect 2448 272 2450 318
rect 2400 210 2450 272
rect 2570 298 2620 340
rect 2570 252 2572 298
rect 2618 252 2620 298
rect 2570 140 2620 252
rect 2740 318 2790 840
rect 2740 272 2742 318
rect 2788 272 2790 318
rect 2740 210 2790 272
rect 0 118 2900 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2900 118
rect 0 0 2900 72
<< via1 >>
rect 104 424 156 476
rect 1304 890 1312 916
rect 1312 890 1356 916
rect 1304 864 1356 890
rect 1634 864 1686 916
rect 374 643 426 646
rect 374 597 377 643
rect 377 597 423 643
rect 423 597 426 643
rect 374 594 426 597
rect 1824 643 1876 646
rect 564 473 616 476
rect 564 427 567 473
rect 567 427 613 473
rect 613 427 616 473
rect 564 424 616 427
rect 944 468 996 476
rect 944 424 947 468
rect 947 424 993 468
rect 993 424 996 468
rect 1824 597 1827 643
rect 1827 597 1873 643
rect 1873 597 1876 643
rect 1824 594 1876 597
rect 1634 513 1686 516
rect 1634 467 1637 513
rect 1637 467 1683 513
rect 1683 467 1686 513
rect 1634 464 1686 467
rect 1304 294 1356 346
rect 1454 334 1506 386
rect 2774 854 2826 906
rect 2614 724 2666 776
rect 2454 583 2506 586
rect 2454 537 2457 583
rect 2457 537 2503 583
rect 2503 537 2506 583
rect 2454 534 2506 537
rect 1894 334 1946 386
rect 2124 354 2176 406
<< metal2 >>
rect 560 1000 1510 1060
rect 350 650 450 660
rect 340 646 460 650
rect 340 594 374 646
rect 426 594 460 646
rect 340 590 460 594
rect 350 580 450 590
rect 560 490 620 1000
rect 1300 930 1360 940
rect 1290 916 1370 930
rect 1290 864 1304 916
rect 1356 864 1370 916
rect 1290 850 1370 864
rect 90 480 170 490
rect 550 480 640 490
rect 930 480 1010 490
rect 80 476 180 480
rect 80 424 104 476
rect 156 424 180 476
rect 80 420 180 424
rect 540 476 640 480
rect 540 424 564 476
rect 616 424 640 476
rect 540 420 640 424
rect 920 476 1020 480
rect 920 424 944 476
rect 996 424 1020 476
rect 920 420 1020 424
rect 90 410 170 420
rect 550 410 640 420
rect 930 410 1010 420
rect 100 290 160 410
rect 940 290 1000 410
rect 1300 360 1360 850
rect 1450 400 1510 1000
rect 1620 920 1700 930
rect 1610 916 2290 920
rect 1610 864 1634 916
rect 1686 864 2290 916
rect 2760 910 2840 920
rect 1610 860 2290 864
rect 1620 850 1700 860
rect 1630 530 1690 850
rect 1810 650 1890 660
rect 1800 646 1900 650
rect 1800 594 1824 646
rect 1876 594 1900 646
rect 1800 590 1900 594
rect 2230 590 2290 860
rect 2750 906 2850 910
rect 2750 854 2774 906
rect 2826 854 2850 906
rect 2750 850 2850 854
rect 2760 840 2840 850
rect 2600 780 2680 790
rect 2590 776 2690 780
rect 2590 724 2614 776
rect 2666 724 2690 776
rect 2590 720 2690 724
rect 2600 710 2680 720
rect 2440 590 2520 600
rect 1810 580 1890 590
rect 2230 586 2530 590
rect 2230 534 2454 586
rect 2506 534 2530 586
rect 2230 530 2530 534
rect 1620 520 1700 530
rect 2440 520 2520 530
rect 1610 516 1710 520
rect 1610 464 1634 516
rect 1686 464 1710 516
rect 1610 460 1710 464
rect 1620 450 1700 460
rect 2110 410 2190 420
rect 2040 406 2200 410
rect 1440 390 1520 400
rect 1880 390 1960 400
rect 1430 386 1980 390
rect 100 230 1000 290
rect 1290 346 1370 360
rect 1290 294 1304 346
rect 1356 294 1370 346
rect 1430 334 1454 386
rect 1506 334 1894 386
rect 1946 334 1980 386
rect 1430 330 1980 334
rect 2040 354 2124 406
rect 2176 354 2200 406
rect 2040 350 2200 354
rect 2040 340 2190 350
rect 1440 320 1520 330
rect 1880 320 1960 330
rect 1290 280 1370 294
rect 1300 260 1370 280
rect 2040 260 2100 340
rect 1300 200 2100 260
<< labels >>
rlabel via1 s 374 594 426 646 4 D
port 1 nsew signal input
rlabel via1 s 2774 854 2826 906 4 Q
port 2 nsew signal output
rlabel via1 s 2614 724 2666 776 4 QN
port 3 nsew signal output
rlabel via1 s 1824 594 1876 646 4 CLK
port 4 nsew clock input
rlabel metal1 s 280 970 330 1270 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 320 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1000 840 1050 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1720 970 1770 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2080 720 2130 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2570 830 2620 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1130 2900 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1000 0 1050 300 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1720 0 1770 320 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2080 0 2130 300 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2570 0 2620 340 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2900 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 1810 580 1890 660 1 CLK
port 4 nsew clock input
rlabel metal2 s 1800 590 1900 650 1 CLK
port 4 nsew clock input
rlabel metal1 s 780 420 840 680 1 CLK
port 4 nsew clock input
rlabel metal1 s 760 420 860 480 1 CLK
port 4 nsew clock input
rlabel metal1 s 1210 410 1270 680 1 CLK
port 4 nsew clock input
rlabel metal1 s 1190 410 1290 470 1 CLK
port 4 nsew clock input
rlabel metal1 s 500 620 1790 680 1 CLK
port 4 nsew clock input
rlabel metal1 s 500 620 1880 670 1 CLK
port 4 nsew clock input
rlabel metal1 s 1800 590 1900 650 1 CLK
port 4 nsew clock input
rlabel metal2 s 350 580 450 660 1 D
port 1 nsew signal input
rlabel metal2 s 340 590 460 650 1 D
port 1 nsew signal input
rlabel metal1 s 350 590 450 650 1 D
port 1 nsew signal input
rlabel metal2 s 2760 840 2840 920 1 Q
port 2 nsew signal output
rlabel metal2 s 2750 850 2850 910 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 210 2790 1060 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 840 2840 920 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 850 2850 920 1 Q
port 2 nsew signal output
rlabel metal2 s 2600 710 2680 790 1 QN
port 3 nsew signal output
rlabel metal2 s 2590 720 2690 780 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 210 2450 440 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 720 2450 1060 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 390 2670 440 1 QN
port 3 nsew signal output
rlabel metal1 s 2610 390 2670 780 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 720 2690 780 1 QN
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2900 1270
string GDS_END 199344
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 178242
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
