magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use nmos_5p0431059130205_512x8m81  nmos_5p0431059130205_512x8m81_0
timestamp 1750858719
transform 1 0 -31 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 256572
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 256322
<< end >>
