magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< metal1 >>
rect 742 2136 1686 2148
rect 742 2084 754 2136
rect 806 2084 878 2136
rect 930 2084 1002 2136
rect 1054 2084 1126 2136
rect 1178 2084 1250 2136
rect 1302 2084 1374 2136
rect 1426 2084 1498 2136
rect 1550 2084 1622 2136
rect 1674 2084 1686 2136
rect 742 2012 1686 2084
rect 742 1960 754 2012
rect 806 1960 878 2012
rect 930 1960 1002 2012
rect 1054 1960 1126 2012
rect 1178 1960 1250 2012
rect 1302 1960 1374 2012
rect 1426 1960 1498 2012
rect 1550 1960 1622 2012
rect 1674 1960 1686 2012
rect 742 1888 1686 1960
rect 742 1836 754 1888
rect 806 1836 878 1888
rect 930 1836 1002 1888
rect 1054 1836 1126 1888
rect 1178 1836 1250 1888
rect 1302 1836 1374 1888
rect 1426 1836 1498 1888
rect 1550 1836 1622 1888
rect 1674 1836 1686 1888
rect 742 1824 1686 1836
<< via1 >>
rect 754 2084 806 2136
rect 878 2084 930 2136
rect 1002 2084 1054 2136
rect 1126 2084 1178 2136
rect 1250 2084 1302 2136
rect 1374 2084 1426 2136
rect 1498 2084 1550 2136
rect 1622 2084 1674 2136
rect 754 1960 806 2012
rect 878 1960 930 2012
rect 1002 1960 1054 2012
rect 1126 1960 1178 2012
rect 1250 1960 1302 2012
rect 1374 1960 1426 2012
rect 1498 1960 1550 2012
rect 1622 1960 1674 2012
rect 754 1836 806 1888
rect 878 1836 930 1888
rect 1002 1836 1054 1888
rect 1126 1836 1178 1888
rect 1250 1836 1302 1888
rect 1374 1836 1426 1888
rect 1498 1836 1550 1888
rect 1622 1836 1674 1888
<< metal2 >>
rect 742 2138 1686 2148
rect 742 2082 752 2138
rect 808 2082 876 2138
rect 932 2082 1000 2138
rect 1056 2082 1124 2138
rect 1180 2082 1248 2138
rect 1304 2082 1372 2138
rect 1428 2082 1496 2138
rect 1552 2082 1620 2138
rect 1676 2082 1686 2138
rect 742 2014 1686 2082
rect 742 1958 752 2014
rect 808 1958 876 2014
rect 932 1958 1000 2014
rect 1056 1958 1124 2014
rect 1180 1958 1248 2014
rect 1304 1958 1372 2014
rect 1428 1958 1496 2014
rect 1552 1958 1620 2014
rect 1676 1958 1686 2014
rect 742 1890 1686 1958
rect 742 1834 752 1890
rect 808 1834 876 1890
rect 932 1834 1000 1890
rect 1056 1834 1124 1890
rect 1180 1834 1248 1890
rect 1304 1834 1372 1890
rect 1428 1834 1496 1890
rect 1552 1834 1620 1890
rect 1676 1834 1686 1890
rect 742 1824 1686 1834
rect -484 1588 460 1598
rect -484 1532 -474 1588
rect -418 1532 -350 1588
rect -294 1532 -226 1588
rect -170 1532 -102 1588
rect -46 1532 22 1588
rect 78 1532 146 1588
rect 202 1532 270 1588
rect 326 1532 394 1588
rect 450 1532 460 1588
rect -484 1464 460 1532
rect -484 1408 -474 1464
rect -418 1408 -350 1464
rect -294 1408 -226 1464
rect -170 1408 -102 1464
rect -46 1408 22 1464
rect 78 1408 146 1464
rect 202 1408 270 1464
rect 326 1408 394 1464
rect 450 1408 460 1464
rect -484 1340 460 1408
rect -484 1284 -474 1340
rect -418 1284 -350 1340
rect -294 1284 -226 1340
rect -170 1284 -102 1340
rect -46 1284 22 1340
rect 78 1284 146 1340
rect 202 1284 270 1340
rect 326 1284 394 1340
rect 450 1284 460 1340
rect -484 1216 460 1284
rect -484 1160 -474 1216
rect -418 1160 -350 1216
rect -294 1160 -226 1216
rect -170 1160 -102 1216
rect -46 1160 22 1216
rect 78 1160 146 1216
rect 202 1160 270 1216
rect 326 1160 394 1216
rect 450 1160 460 1216
rect -484 1092 460 1160
rect -484 1036 -474 1092
rect -418 1036 -350 1092
rect -294 1036 -226 1092
rect -170 1036 -102 1092
rect -46 1036 22 1092
rect 78 1036 146 1092
rect 202 1036 270 1092
rect 326 1036 394 1092
rect 450 1036 460 1092
rect -484 968 460 1036
rect -484 912 -474 968
rect -418 912 -350 968
rect -294 912 -226 968
rect -170 912 -102 968
rect -46 912 22 968
rect 78 912 146 968
rect 202 912 270 968
rect 326 912 394 968
rect 450 912 460 968
rect -484 844 460 912
rect -484 788 -474 844
rect -418 788 -350 844
rect -294 788 -226 844
rect -170 788 -102 844
rect -46 788 22 844
rect 78 788 146 844
rect 202 788 270 844
rect 326 788 394 844
rect 450 788 460 844
rect -484 720 460 788
rect -484 664 -474 720
rect -418 664 -350 720
rect -294 664 -226 720
rect -170 664 -102 720
rect -46 664 22 720
rect 78 664 146 720
rect 202 664 270 720
rect 326 664 394 720
rect 450 664 460 720
rect -484 654 460 664
<< via2 >>
rect 752 2136 808 2138
rect 752 2084 754 2136
rect 754 2084 806 2136
rect 806 2084 808 2136
rect 752 2082 808 2084
rect 876 2136 932 2138
rect 876 2084 878 2136
rect 878 2084 930 2136
rect 930 2084 932 2136
rect 876 2082 932 2084
rect 1000 2136 1056 2138
rect 1000 2084 1002 2136
rect 1002 2084 1054 2136
rect 1054 2084 1056 2136
rect 1000 2082 1056 2084
rect 1124 2136 1180 2138
rect 1124 2084 1126 2136
rect 1126 2084 1178 2136
rect 1178 2084 1180 2136
rect 1124 2082 1180 2084
rect 1248 2136 1304 2138
rect 1248 2084 1250 2136
rect 1250 2084 1302 2136
rect 1302 2084 1304 2136
rect 1248 2082 1304 2084
rect 1372 2136 1428 2138
rect 1372 2084 1374 2136
rect 1374 2084 1426 2136
rect 1426 2084 1428 2136
rect 1372 2082 1428 2084
rect 1496 2136 1552 2138
rect 1496 2084 1498 2136
rect 1498 2084 1550 2136
rect 1550 2084 1552 2136
rect 1496 2082 1552 2084
rect 1620 2136 1676 2138
rect 1620 2084 1622 2136
rect 1622 2084 1674 2136
rect 1674 2084 1676 2136
rect 1620 2082 1676 2084
rect 752 2012 808 2014
rect 752 1960 754 2012
rect 754 1960 806 2012
rect 806 1960 808 2012
rect 752 1958 808 1960
rect 876 2012 932 2014
rect 876 1960 878 2012
rect 878 1960 930 2012
rect 930 1960 932 2012
rect 876 1958 932 1960
rect 1000 2012 1056 2014
rect 1000 1960 1002 2012
rect 1002 1960 1054 2012
rect 1054 1960 1056 2012
rect 1000 1958 1056 1960
rect 1124 2012 1180 2014
rect 1124 1960 1126 2012
rect 1126 1960 1178 2012
rect 1178 1960 1180 2012
rect 1124 1958 1180 1960
rect 1248 2012 1304 2014
rect 1248 1960 1250 2012
rect 1250 1960 1302 2012
rect 1302 1960 1304 2012
rect 1248 1958 1304 1960
rect 1372 2012 1428 2014
rect 1372 1960 1374 2012
rect 1374 1960 1426 2012
rect 1426 1960 1428 2012
rect 1372 1958 1428 1960
rect 1496 2012 1552 2014
rect 1496 1960 1498 2012
rect 1498 1960 1550 2012
rect 1550 1960 1552 2012
rect 1496 1958 1552 1960
rect 1620 2012 1676 2014
rect 1620 1960 1622 2012
rect 1622 1960 1674 2012
rect 1674 1960 1676 2012
rect 1620 1958 1676 1960
rect 752 1888 808 1890
rect 752 1836 754 1888
rect 754 1836 806 1888
rect 806 1836 808 1888
rect 752 1834 808 1836
rect 876 1888 932 1890
rect 876 1836 878 1888
rect 878 1836 930 1888
rect 930 1836 932 1888
rect 876 1834 932 1836
rect 1000 1888 1056 1890
rect 1000 1836 1002 1888
rect 1002 1836 1054 1888
rect 1054 1836 1056 1888
rect 1000 1834 1056 1836
rect 1124 1888 1180 1890
rect 1124 1836 1126 1888
rect 1126 1836 1178 1888
rect 1178 1836 1180 1888
rect 1124 1834 1180 1836
rect 1248 1888 1304 1890
rect 1248 1836 1250 1888
rect 1250 1836 1302 1888
rect 1302 1836 1304 1888
rect 1248 1834 1304 1836
rect 1372 1888 1428 1890
rect 1372 1836 1374 1888
rect 1374 1836 1426 1888
rect 1426 1836 1428 1888
rect 1372 1834 1428 1836
rect 1496 1888 1552 1890
rect 1496 1836 1498 1888
rect 1498 1836 1550 1888
rect 1550 1836 1552 1888
rect 1496 1834 1552 1836
rect 1620 1888 1676 1890
rect 1620 1836 1622 1888
rect 1622 1836 1674 1888
rect 1674 1836 1676 1888
rect 1620 1834 1676 1836
rect -474 1532 -418 1588
rect -350 1532 -294 1588
rect -226 1532 -170 1588
rect -102 1532 -46 1588
rect 22 1532 78 1588
rect 146 1532 202 1588
rect 270 1532 326 1588
rect 394 1532 450 1588
rect -474 1408 -418 1464
rect -350 1408 -294 1464
rect -226 1408 -170 1464
rect -102 1408 -46 1464
rect 22 1408 78 1464
rect 146 1408 202 1464
rect 270 1408 326 1464
rect 394 1408 450 1464
rect -474 1284 -418 1340
rect -350 1284 -294 1340
rect -226 1284 -170 1340
rect -102 1284 -46 1340
rect 22 1284 78 1340
rect 146 1284 202 1340
rect 270 1284 326 1340
rect 394 1284 450 1340
rect -474 1160 -418 1216
rect -350 1160 -294 1216
rect -226 1160 -170 1216
rect -102 1160 -46 1216
rect 22 1160 78 1216
rect 146 1160 202 1216
rect 270 1160 326 1216
rect 394 1160 450 1216
rect -474 1036 -418 1092
rect -350 1036 -294 1092
rect -226 1036 -170 1092
rect -102 1036 -46 1092
rect 22 1036 78 1092
rect 146 1036 202 1092
rect 270 1036 326 1092
rect 394 1036 450 1092
rect -474 912 -418 968
rect -350 912 -294 968
rect -226 912 -170 968
rect -102 912 -46 968
rect 22 912 78 968
rect 146 912 202 968
rect 270 912 326 968
rect 394 912 450 968
rect -474 788 -418 844
rect -350 788 -294 844
rect -226 788 -170 844
rect -102 788 -46 844
rect 22 788 78 844
rect 146 788 202 844
rect 270 788 326 844
rect 394 788 450 844
rect -474 664 -418 720
rect -350 664 -294 720
rect -226 664 -170 720
rect -102 664 -46 720
rect 22 664 78 720
rect 146 664 202 720
rect 270 664 326 720
rect 394 664 450 720
<< metal3 >>
rect -511 1588 489 2430
rect 714 2138 1714 2430
rect 714 2082 752 2138
rect 808 2082 876 2138
rect 932 2082 1000 2138
rect 1056 2082 1124 2138
rect 1180 2082 1248 2138
rect 1304 2082 1372 2138
rect 1428 2082 1496 2138
rect 1552 2082 1620 2138
rect 1676 2082 1714 2138
rect 714 2014 1714 2082
rect 714 1958 752 2014
rect 808 1958 876 2014
rect 932 1958 1000 2014
rect 1056 1958 1124 2014
rect 1180 1958 1248 2014
rect 1304 1958 1372 2014
rect 1428 1958 1496 2014
rect 1552 1958 1620 2014
rect 1676 1958 1714 2014
rect 714 1890 1714 1958
rect 714 1834 752 1890
rect 808 1834 876 1890
rect 932 1834 1000 1890
rect 1056 1834 1124 1890
rect 1180 1834 1248 1890
rect 1304 1834 1372 1890
rect 1428 1834 1496 1890
rect 1552 1834 1620 1890
rect 1676 1834 1714 1890
rect 714 1822 1714 1834
rect -511 1532 -474 1588
rect -418 1532 -350 1588
rect -294 1532 -226 1588
rect -170 1532 -102 1588
rect -46 1532 22 1588
rect 78 1532 146 1588
rect 202 1532 270 1588
rect 326 1532 394 1588
rect 450 1532 489 1588
rect -511 1464 489 1532
rect -511 1408 -474 1464
rect -418 1408 -350 1464
rect -294 1408 -226 1464
rect -170 1408 -102 1464
rect -46 1408 22 1464
rect 78 1408 146 1464
rect 202 1408 270 1464
rect 326 1408 394 1464
rect 450 1408 489 1464
rect -511 1340 489 1408
rect -511 1284 -474 1340
rect -418 1284 -350 1340
rect -294 1284 -226 1340
rect -170 1284 -102 1340
rect -46 1284 22 1340
rect 78 1284 146 1340
rect 202 1284 270 1340
rect 326 1284 394 1340
rect 450 1284 489 1340
rect -511 1216 489 1284
rect -511 1160 -474 1216
rect -418 1160 -350 1216
rect -294 1160 -226 1216
rect -170 1160 -102 1216
rect -46 1160 22 1216
rect 78 1160 146 1216
rect 202 1160 270 1216
rect 326 1160 394 1216
rect 450 1160 489 1216
rect -511 1092 489 1160
rect -511 1036 -474 1092
rect -418 1036 -350 1092
rect -294 1036 -226 1092
rect -170 1036 -102 1092
rect -46 1036 22 1092
rect 78 1036 146 1092
rect 202 1036 270 1092
rect 326 1036 394 1092
rect 450 1036 489 1092
rect -511 968 489 1036
rect -511 912 -474 968
rect -418 912 -350 968
rect -294 912 -226 968
rect -170 912 -102 968
rect -46 912 22 968
rect 78 912 146 968
rect 202 912 270 968
rect 326 912 394 968
rect 450 912 489 968
rect -511 844 489 912
rect -511 788 -474 844
rect -418 788 -350 844
rect -294 788 -226 844
rect -170 788 -102 844
rect -46 788 22 844
rect 78 788 146 844
rect 202 788 270 844
rect 326 788 394 844
rect 450 788 489 844
rect -511 720 489 788
rect -511 664 -474 720
rect -418 664 -350 720
rect -294 664 -226 720
rect -170 664 -102 720
rect -46 664 22 720
rect 78 664 146 720
rect 202 664 270 720
rect 326 664 394 720
rect 450 664 489 720
rect -511 630 489 664
use M2_M14310590878179_256x8m81  M2_M14310590878179_256x8m81_0
timestamp 1750858719
transform 1 0 1214 0 1 1986
box 0 0 1 1
use M3_M24310590878178_256x8m81  M3_M24310590878178_256x8m81_0
timestamp 1750858719
transform 1 0 1214 0 1 1986
box 0 0 1 1
use M3_M24310590878180_256x8m81  M3_M24310590878180_256x8m81_0
timestamp 1750858719
transform 1 0 -12 0 1 1126
box 0 0 1 1
<< properties >>
string GDS_END 2396384
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2396116
string path -0.055 3.150 -0.055 12.150 
<< end >>
