magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 377 1766 870
rect -86 352 882 377
rect 1139 352 1766 377
<< pwell >>
rect -86 -86 1766 352
<< metal1 >>
rect 0 724 1680 844
rect 49 506 95 724
rect 141 305 200 664
rect 360 305 424 664
rect 584 305 648 664
rect 49 60 95 163
rect 497 60 543 163
rect 698 244 758 676
rect 808 305 872 664
rect 1032 428 1096 664
rect 1256 428 1320 664
rect 1461 506 1507 724
rect 1032 354 1208 428
rect 1256 354 1574 428
rect 698 198 1527 244
rect 1481 111 1527 198
rect 0 -60 1680 60
<< obsm1 >>
rect 273 209 635 255
rect 273 106 319 209
rect 589 152 635 209
rect 589 106 1314 152
<< labels >>
rlabel metal1 s 808 305 872 664 6 A1
port 1 nsew default input
rlabel metal1 s 1032 354 1208 428 6 A2
port 2 nsew default input
rlabel metal1 s 1032 428 1096 664 6 A2
port 2 nsew default input
rlabel metal1 s 1256 354 1574 428 6 A3
port 3 nsew default input
rlabel metal1 s 1256 428 1320 664 6 A3
port 3 nsew default input
rlabel metal1 s 584 305 648 664 6 B1
port 4 nsew default input
rlabel metal1 s 360 305 424 664 6 B2
port 5 nsew default input
rlabel metal1 s 141 305 200 664 6 B3
port 6 nsew default input
rlabel metal1 s 1481 111 1527 198 6 ZN
port 7 nsew default output
rlabel metal1 s 698 198 1527 244 6 ZN
port 7 nsew default output
rlabel metal1 s 698 244 758 676 6 ZN
port 7 nsew default output
rlabel metal1 s 1461 506 1507 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 724 1680 844 6 VDD
port 8 nsew power bidirectional abutment
rlabel nwell s 1139 352 1766 377 6 VNW
port 9 nsew power bidirectional
rlabel nwell s -86 352 882 377 6 VNW
port 9 nsew power bidirectional
rlabel nwell s -86 377 1766 870 6 VNW
port 9 nsew power bidirectional
rlabel pwell s -86 -86 1766 352 6 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 0 -60 1680 60 8 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 163 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 163 6 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1680 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 73490
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 69256
<< end >>
