magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 407 6582 870
rect -86 352 575 407
rect 949 352 6582 407
<< pwell >>
rect 575 352 949 407
rect -86 -86 6582 352
<< mvnmos >>
rect 124 69 244 232
rect 348 69 468 232
rect 572 69 692 232
rect 1064 68 1184 232
rect 1288 68 1408 232
rect 1512 68 1632 232
rect 1736 68 1856 232
rect 1960 68 2080 232
rect 2184 68 2304 232
rect 2408 68 2528 232
rect 2632 68 2752 232
rect 2856 68 2976 232
rect 3080 68 3200 232
rect 3304 68 3424 232
rect 3528 68 3648 232
rect 3752 68 3872 232
rect 3976 68 4096 232
rect 4200 68 4320 232
rect 4424 68 4544 232
rect 4648 68 4768 232
rect 4872 68 4992 232
rect 5096 68 5216 232
rect 5320 68 5440 232
rect 5544 68 5664 232
rect 5768 68 5888 232
rect 5992 68 6112 232
rect 6216 68 6336 232
<< mvpmos >>
rect 172 527 272 711
rect 376 527 476 711
rect 660 527 760 711
rect 1144 481 1244 711
rect 1348 481 1448 711
rect 1552 481 1652 711
rect 1756 481 1856 711
rect 1960 481 2060 711
rect 2224 481 2324 711
rect 2428 481 2528 711
rect 2668 481 2768 716
rect 2872 481 2972 716
rect 3076 481 3176 716
rect 3280 481 3380 716
rect 3484 481 3584 716
rect 3688 481 3788 716
rect 3892 481 3992 716
rect 4096 481 4196 716
rect 4300 481 4400 716
rect 4504 481 4604 716
rect 4708 481 4808 716
rect 4912 481 5012 716
rect 5116 481 5216 716
rect 5320 481 5420 716
rect 5524 481 5624 716
rect 5728 481 5828 716
rect 5932 481 6032 716
<< mvndiff >>
rect 752 274 824 287
rect 752 232 765 274
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 69 124 173
rect 244 128 348 232
rect 244 82 273 128
rect 319 82 348 128
rect 244 69 348 82
rect 468 169 572 232
rect 468 123 497 169
rect 543 123 572 169
rect 468 69 572 123
rect 692 228 765 232
rect 811 228 824 274
rect 692 69 824 228
rect 932 95 1064 232
rect 932 49 945 95
rect 991 68 1064 95
rect 1184 219 1288 232
rect 1184 173 1213 219
rect 1259 173 1288 219
rect 1184 68 1288 173
rect 1408 127 1512 232
rect 1408 81 1437 127
rect 1483 81 1512 127
rect 1408 68 1512 81
rect 1632 219 1736 232
rect 1632 173 1661 219
rect 1707 173 1736 219
rect 1632 68 1736 173
rect 1856 127 1960 232
rect 1856 81 1885 127
rect 1931 81 1960 127
rect 1856 68 1960 81
rect 2080 219 2184 232
rect 2080 173 2109 219
rect 2155 173 2184 219
rect 2080 68 2184 173
rect 2304 127 2408 232
rect 2304 81 2333 127
rect 2379 81 2408 127
rect 2304 68 2408 81
rect 2528 219 2632 232
rect 2528 173 2557 219
rect 2603 173 2632 219
rect 2528 68 2632 173
rect 2752 127 2856 232
rect 2752 81 2781 127
rect 2827 81 2856 127
rect 2752 68 2856 81
rect 2976 219 3080 232
rect 2976 173 3005 219
rect 3051 173 3080 219
rect 2976 68 3080 173
rect 3200 127 3304 232
rect 3200 81 3229 127
rect 3275 81 3304 127
rect 3200 68 3304 81
rect 3424 219 3528 232
rect 3424 173 3453 219
rect 3499 173 3528 219
rect 3424 68 3528 173
rect 3648 127 3752 232
rect 3648 81 3677 127
rect 3723 81 3752 127
rect 3648 68 3752 81
rect 3872 219 3976 232
rect 3872 173 3901 219
rect 3947 173 3976 219
rect 3872 68 3976 173
rect 4096 127 4200 232
rect 4096 81 4125 127
rect 4171 81 4200 127
rect 4096 68 4200 81
rect 4320 219 4424 232
rect 4320 173 4349 219
rect 4395 173 4424 219
rect 4320 68 4424 173
rect 4544 127 4648 232
rect 4544 81 4573 127
rect 4619 81 4648 127
rect 4544 68 4648 81
rect 4768 219 4872 232
rect 4768 173 4797 219
rect 4843 173 4872 219
rect 4768 68 4872 173
rect 4992 127 5096 232
rect 4992 81 5021 127
rect 5067 81 5096 127
rect 4992 68 5096 81
rect 5216 219 5320 232
rect 5216 173 5245 219
rect 5291 173 5320 219
rect 5216 68 5320 173
rect 5440 127 5544 232
rect 5440 81 5469 127
rect 5515 81 5544 127
rect 5440 68 5544 81
rect 5664 219 5768 232
rect 5664 173 5693 219
rect 5739 173 5768 219
rect 5664 68 5768 173
rect 5888 127 5992 232
rect 5888 81 5917 127
rect 5963 81 5992 127
rect 5888 68 5992 81
rect 6112 219 6216 232
rect 6112 173 6141 219
rect 6187 173 6216 219
rect 6112 68 6216 173
rect 6336 141 6424 232
rect 6336 95 6365 141
rect 6411 95 6424 141
rect 6336 68 6424 95
rect 991 49 1004 68
rect 932 36 1004 49
<< mvpdiff >>
rect 2588 711 2668 716
rect 84 602 172 711
rect 84 556 97 602
rect 143 556 172 602
rect 84 527 172 556
rect 272 698 376 711
rect 272 652 301 698
rect 347 652 376 698
rect 272 527 376 652
rect 476 678 660 711
rect 476 632 557 678
rect 603 632 660 678
rect 476 527 660 632
rect 760 586 848 711
rect 760 540 789 586
rect 835 540 848 586
rect 760 527 848 540
rect 1056 665 1144 711
rect 1056 619 1069 665
rect 1115 619 1144 665
rect 1056 481 1144 619
rect 1244 665 1348 711
rect 1244 525 1273 665
rect 1319 525 1348 665
rect 1244 481 1348 525
rect 1448 665 1552 711
rect 1448 619 1477 665
rect 1523 619 1552 665
rect 1448 481 1552 619
rect 1652 665 1756 711
rect 1652 525 1681 665
rect 1727 525 1756 665
rect 1652 481 1756 525
rect 1856 665 1960 711
rect 1856 619 1885 665
rect 1931 619 1960 665
rect 1856 481 1960 619
rect 2060 665 2224 711
rect 2060 525 2120 665
rect 2166 525 2224 665
rect 2060 481 2224 525
rect 2324 665 2428 711
rect 2324 619 2353 665
rect 2399 619 2428 665
rect 2324 481 2428 619
rect 2528 665 2668 711
rect 2528 525 2569 665
rect 2615 525 2668 665
rect 2528 481 2668 525
rect 2768 665 2872 716
rect 2768 525 2797 665
rect 2843 525 2872 665
rect 2768 481 2872 525
rect 2972 665 3076 716
rect 2972 525 3001 665
rect 3047 525 3076 665
rect 2972 481 3076 525
rect 3176 703 3280 716
rect 3176 657 3205 703
rect 3251 657 3280 703
rect 3176 481 3280 657
rect 3380 665 3484 716
rect 3380 525 3409 665
rect 3455 525 3484 665
rect 3380 481 3484 525
rect 3584 703 3688 716
rect 3584 657 3613 703
rect 3659 657 3688 703
rect 3584 481 3688 657
rect 3788 665 3892 716
rect 3788 525 3817 665
rect 3863 525 3892 665
rect 3788 481 3892 525
rect 3992 703 4096 716
rect 3992 657 4021 703
rect 4067 657 4096 703
rect 3992 481 4096 657
rect 4196 665 4300 716
rect 4196 525 4225 665
rect 4271 525 4300 665
rect 4196 481 4300 525
rect 4400 703 4504 716
rect 4400 657 4429 703
rect 4475 657 4504 703
rect 4400 481 4504 657
rect 4604 665 4708 716
rect 4604 525 4633 665
rect 4679 525 4708 665
rect 4604 481 4708 525
rect 4808 703 4912 716
rect 4808 657 4837 703
rect 4883 657 4912 703
rect 4808 481 4912 657
rect 5012 665 5116 716
rect 5012 525 5041 665
rect 5087 525 5116 665
rect 5012 481 5116 525
rect 5216 703 5320 716
rect 5216 657 5245 703
rect 5291 657 5320 703
rect 5216 481 5320 657
rect 5420 665 5524 716
rect 5420 525 5449 665
rect 5495 525 5524 665
rect 5420 481 5524 525
rect 5624 703 5728 716
rect 5624 657 5653 703
rect 5699 657 5728 703
rect 5624 481 5728 657
rect 5828 665 5932 716
rect 5828 525 5857 665
rect 5903 525 5932 665
rect 5828 481 5932 525
rect 6032 665 6120 716
rect 6032 525 6061 665
rect 6107 525 6120 665
rect 6032 481 6120 525
<< mvndiffc >>
rect 49 173 95 219
rect 273 82 319 128
rect 497 123 543 169
rect 765 228 811 274
rect 945 49 991 95
rect 1213 173 1259 219
rect 1437 81 1483 127
rect 1661 173 1707 219
rect 1885 81 1931 127
rect 2109 173 2155 219
rect 2333 81 2379 127
rect 2557 173 2603 219
rect 2781 81 2827 127
rect 3005 173 3051 219
rect 3229 81 3275 127
rect 3453 173 3499 219
rect 3677 81 3723 127
rect 3901 173 3947 219
rect 4125 81 4171 127
rect 4349 173 4395 219
rect 4573 81 4619 127
rect 4797 173 4843 219
rect 5021 81 5067 127
rect 5245 173 5291 219
rect 5469 81 5515 127
rect 5693 173 5739 219
rect 5917 81 5963 127
rect 6141 173 6187 219
rect 6365 95 6411 141
<< mvpdiffc >>
rect 97 556 143 602
rect 301 652 347 698
rect 557 632 603 678
rect 789 540 835 586
rect 1069 619 1115 665
rect 1273 525 1319 665
rect 1477 619 1523 665
rect 1681 525 1727 665
rect 1885 619 1931 665
rect 2120 525 2166 665
rect 2353 619 2399 665
rect 2569 525 2615 665
rect 2797 525 2843 665
rect 3001 525 3047 665
rect 3205 657 3251 703
rect 3409 525 3455 665
rect 3613 657 3659 703
rect 3817 525 3863 665
rect 4021 657 4067 703
rect 4225 525 4271 665
rect 4429 657 4475 703
rect 4633 525 4679 665
rect 4837 657 4883 703
rect 5041 525 5087 665
rect 5245 657 5291 703
rect 5449 525 5495 665
rect 5653 657 5699 703
rect 5857 525 5903 665
rect 6061 525 6107 665
<< polysilicon >>
rect 172 711 272 755
rect 376 711 476 755
rect 660 711 760 755
rect 1144 711 1244 755
rect 1348 711 1448 755
rect 1552 711 1652 755
rect 1756 711 1856 755
rect 1960 711 2060 755
rect 2224 711 2324 755
rect 2428 711 2528 755
rect 2668 716 2768 760
rect 2872 716 2972 760
rect 3076 716 3176 760
rect 3280 716 3380 760
rect 3484 716 3584 760
rect 3688 716 3788 760
rect 3892 716 3992 760
rect 4096 716 4196 760
rect 4300 716 4400 760
rect 4504 716 4604 760
rect 4708 716 4808 760
rect 4912 716 5012 760
rect 5116 716 5216 760
rect 5320 716 5420 760
rect 5524 716 5624 760
rect 5728 716 5828 760
rect 5932 716 6032 760
rect 172 413 272 527
rect 376 413 476 527
rect 660 493 760 527
rect 660 447 673 493
rect 719 447 760 493
rect 660 434 760 447
rect 172 412 612 413
rect 172 366 185 412
rect 231 373 612 412
rect 231 366 244 373
rect 172 288 244 366
rect 124 232 244 288
rect 348 311 468 324
rect 348 265 379 311
rect 425 265 468 311
rect 348 232 468 265
rect 572 288 612 373
rect 1144 401 1244 481
rect 1144 355 1171 401
rect 1217 363 1244 401
rect 1348 401 1448 481
rect 1348 363 1373 401
rect 1217 355 1373 363
rect 1419 363 1448 401
rect 1552 401 1652 481
rect 1552 363 1578 401
rect 1419 355 1578 363
rect 1624 363 1652 401
rect 1756 401 1856 481
rect 1756 363 1781 401
rect 1624 355 1781 363
rect 1827 363 1856 401
rect 1960 401 2060 481
rect 1960 363 1987 401
rect 1827 355 1987 363
rect 2033 363 2060 401
rect 2224 401 2324 481
rect 2224 363 2251 401
rect 2033 355 2251 363
rect 2297 363 2324 401
rect 2428 401 2528 481
rect 2428 363 2455 401
rect 2297 355 2455 363
rect 2501 363 2528 401
rect 2668 363 2768 481
rect 2872 446 2972 481
rect 2872 400 2902 446
rect 2948 420 2972 446
rect 3076 446 3176 481
rect 3076 420 3105 446
rect 2948 400 3105 420
rect 3151 420 3176 446
rect 3280 446 3380 481
rect 3280 420 3309 446
rect 3151 400 3309 420
rect 3355 420 3380 446
rect 3484 446 3584 481
rect 3484 420 3513 446
rect 3355 400 3513 420
rect 3559 420 3584 446
rect 3688 446 3788 481
rect 3688 420 3715 446
rect 3559 400 3715 420
rect 3761 420 3788 446
rect 3892 446 3992 481
rect 3892 420 3919 446
rect 3761 400 3919 420
rect 3965 420 3992 446
rect 4096 446 4196 481
rect 4096 420 4124 446
rect 3965 400 4124 420
rect 4170 420 4196 446
rect 4300 446 4400 481
rect 4300 420 4327 446
rect 4170 400 4327 420
rect 4373 420 4400 446
rect 4504 420 4604 481
rect 4708 446 4808 481
rect 4708 420 4737 446
rect 4373 400 4737 420
rect 4783 420 4808 446
rect 4912 446 5012 481
rect 4912 420 4940 446
rect 4783 400 4940 420
rect 4986 420 5012 446
rect 5116 446 5216 481
rect 5116 420 5144 446
rect 4986 400 5144 420
rect 5190 420 5216 446
rect 5320 446 5420 481
rect 5320 420 5346 446
rect 5190 400 5346 420
rect 5392 420 5420 446
rect 5524 446 5624 481
rect 5524 420 5553 446
rect 5392 400 5553 420
rect 5599 420 5624 446
rect 5728 446 5828 481
rect 5728 420 5752 446
rect 5599 400 5752 420
rect 5798 420 5828 446
rect 5932 446 6032 481
rect 5932 420 5959 446
rect 5798 400 5959 420
rect 6005 400 6032 446
rect 2872 380 6032 400
rect 2501 355 2768 363
rect 1144 342 2768 355
rect 1144 323 2752 342
rect 572 232 692 288
rect 1144 287 1184 323
rect 1064 232 1184 287
rect 1288 232 1408 323
rect 1512 232 1632 323
rect 1736 232 1856 323
rect 1960 232 2080 323
rect 2184 232 2304 323
rect 2408 232 2528 323
rect 2632 232 2752 323
rect 2856 318 6336 332
rect 2856 272 2869 318
rect 2915 292 3118 318
rect 2915 272 2976 292
rect 2856 232 2976 272
rect 3080 272 3118 292
rect 3164 292 3341 318
rect 3164 272 3200 292
rect 3080 232 3200 272
rect 3304 272 3341 292
rect 3387 292 3564 318
rect 3387 272 3424 292
rect 3304 232 3424 272
rect 3528 272 3564 292
rect 3610 292 3789 318
rect 3610 272 3648 292
rect 3528 232 3648 272
rect 3752 272 3789 292
rect 3835 292 4014 318
rect 3835 272 3872 292
rect 3752 232 3872 272
rect 3976 272 4014 292
rect 4060 292 4233 318
rect 4060 272 4096 292
rect 3976 232 4096 272
rect 4200 272 4233 292
rect 4279 292 4709 318
rect 4279 272 4320 292
rect 4200 232 4320 272
rect 4424 232 4544 292
rect 4648 272 4709 292
rect 4755 292 4910 318
rect 4755 272 4768 292
rect 4648 232 4768 272
rect 4872 272 4910 292
rect 4956 292 5134 318
rect 4956 272 4992 292
rect 4872 232 4992 272
rect 5096 272 5134 292
rect 5180 292 5356 318
rect 5180 272 5216 292
rect 5096 232 5216 272
rect 5320 272 5356 292
rect 5402 292 5584 318
rect 5402 272 5440 292
rect 5320 232 5440 272
rect 5544 272 5584 292
rect 5630 292 5797 318
rect 5630 272 5664 292
rect 5544 232 5664 272
rect 5768 272 5797 292
rect 5843 292 6019 318
rect 5843 272 5888 292
rect 5768 232 5888 272
rect 5992 272 6019 292
rect 6065 292 6247 318
rect 6065 272 6112 292
rect 5992 232 6112 272
rect 6216 272 6247 292
rect 6293 272 6336 318
rect 6216 232 6336 272
rect 124 24 244 69
rect 348 24 468 69
rect 572 24 692 69
rect 1064 24 1184 68
rect 1288 24 1408 68
rect 1512 24 1632 68
rect 1736 24 1856 68
rect 1960 24 2080 68
rect 2184 24 2304 68
rect 2408 24 2528 68
rect 2632 24 2752 68
rect 2856 24 2976 68
rect 3080 24 3200 68
rect 3304 24 3424 68
rect 3528 24 3648 68
rect 3752 24 3872 68
rect 3976 24 4096 68
rect 4200 24 4320 68
rect 4424 24 4544 68
rect 4648 24 4768 68
rect 4872 24 4992 68
rect 5096 24 5216 68
rect 5320 24 5440 68
rect 5544 24 5664 68
rect 5768 24 5888 68
rect 5992 24 6112 68
rect 6216 24 6336 68
<< polycontact >>
rect 673 447 719 493
rect 185 366 231 412
rect 379 265 425 311
rect 1171 355 1217 401
rect 1373 355 1419 401
rect 1578 355 1624 401
rect 1781 355 1827 401
rect 1987 355 2033 401
rect 2251 355 2297 401
rect 2455 355 2501 401
rect 2902 400 2948 446
rect 3105 400 3151 446
rect 3309 400 3355 446
rect 3513 400 3559 446
rect 3715 400 3761 446
rect 3919 400 3965 446
rect 4124 400 4170 446
rect 4327 400 4373 446
rect 4737 400 4783 446
rect 4940 400 4986 446
rect 5144 400 5190 446
rect 5346 400 5392 446
rect 5553 400 5599 446
rect 5752 400 5798 446
rect 5959 400 6005 446
rect 2869 272 2915 318
rect 3118 272 3164 318
rect 3341 272 3387 318
rect 3564 272 3610 318
rect 3789 272 3835 318
rect 4014 272 4060 318
rect 4233 272 4279 318
rect 4709 272 4755 318
rect 4910 272 4956 318
rect 5134 272 5180 318
rect 5356 272 5402 318
rect 5584 272 5630 318
rect 5797 272 5843 318
rect 6019 272 6065 318
rect 6247 272 6293 318
<< metal1 >>
rect 0 724 6496 844
rect 290 698 358 724
rect 290 652 301 698
rect 347 652 358 698
rect 546 632 557 678
rect 603 632 1012 678
rect 84 556 97 602
rect 143 556 425 602
rect 379 504 425 556
rect 778 540 789 586
rect 835 540 846 586
rect 379 493 730 504
rect 379 447 673 493
rect 719 447 730 493
rect 74 412 318 430
rect 74 366 185 412
rect 231 366 318 412
rect 74 354 318 366
rect 379 311 425 447
rect 778 401 846 540
rect 38 219 425 265
rect 497 355 846 401
rect 966 552 1012 632
rect 1058 665 1126 724
rect 1058 619 1069 665
rect 1115 619 1126 665
rect 1058 608 1126 619
rect 1262 665 1330 676
rect 1262 552 1273 665
rect 966 525 1273 552
rect 1319 552 1330 665
rect 1466 665 1534 724
rect 1466 619 1477 665
rect 1523 619 1534 665
rect 1466 608 1534 619
rect 1670 665 1738 676
rect 1670 552 1681 665
rect 1319 525 1681 552
rect 1727 552 1738 665
rect 1874 665 1942 724
rect 1874 619 1885 665
rect 1931 619 1942 665
rect 1874 608 1942 619
rect 2109 665 2177 676
rect 2109 552 2120 665
rect 1727 525 2120 552
rect 2166 552 2177 665
rect 2342 665 2410 724
rect 2342 619 2353 665
rect 2399 619 2410 665
rect 2342 608 2410 619
rect 2558 665 2626 676
rect 2558 552 2569 665
rect 2166 525 2569 552
rect 2615 552 2626 665
rect 2786 665 2854 724
rect 3194 703 3262 724
rect 2615 525 2723 552
rect 966 506 2723 525
rect 2786 525 2797 665
rect 2843 525 2854 665
rect 2786 506 2854 525
rect 2990 665 3058 676
rect 2990 525 3001 665
rect 3047 611 3058 665
rect 3194 657 3205 703
rect 3251 657 3262 703
rect 3602 703 3670 724
rect 3398 665 3466 676
rect 3398 611 3409 665
rect 3047 525 3409 611
rect 3455 611 3466 665
rect 3602 657 3613 703
rect 3659 657 3670 703
rect 4010 703 4078 724
rect 3806 665 3874 676
rect 3806 611 3817 665
rect 3455 525 3817 611
rect 3863 611 3874 665
rect 4010 657 4021 703
rect 4067 657 4078 703
rect 4418 703 4486 724
rect 4214 665 4282 676
rect 4214 611 4225 665
rect 3863 525 4225 611
rect 4271 611 4282 665
rect 4418 657 4429 703
rect 4475 657 4486 703
rect 4826 703 4894 724
rect 4626 665 4690 676
rect 4626 611 4633 665
rect 4271 525 4633 611
rect 4679 611 4690 665
rect 4826 657 4837 703
rect 4883 657 4894 703
rect 5234 703 5302 724
rect 5030 665 5098 676
rect 5030 611 5041 665
rect 4679 525 5041 611
rect 5087 611 5098 665
rect 5234 657 5245 703
rect 5291 657 5302 703
rect 5642 703 5710 724
rect 5438 665 5506 676
rect 5438 611 5449 665
rect 5087 525 5449 611
rect 5495 611 5506 665
rect 5642 657 5653 703
rect 5699 657 5710 703
rect 5846 665 5914 676
rect 5846 611 5857 665
rect 5495 525 5857 611
rect 5903 525 5914 665
rect 38 173 49 219
rect 95 173 106 219
rect 497 169 543 355
rect 966 309 1012 506
rect 2654 446 2723 506
rect 2990 501 5914 525
rect 6061 665 6107 724
rect 6061 506 6107 525
rect 1138 401 2558 430
rect 1138 355 1171 401
rect 1217 355 1373 401
rect 1419 355 1578 401
rect 1624 355 1781 401
rect 1827 355 1987 401
rect 2033 355 2251 401
rect 2297 355 2455 401
rect 2501 355 2558 401
rect 2654 400 2902 446
rect 2948 400 3105 446
rect 3151 400 3309 446
rect 3355 400 3513 446
rect 3559 400 3715 446
rect 3761 400 3919 446
rect 3965 400 4124 446
rect 4170 400 4327 446
rect 4373 400 4384 446
rect 1138 354 2558 355
rect 754 274 1012 309
rect 754 228 765 274
rect 811 263 1012 274
rect 2670 272 2869 318
rect 2915 272 3118 318
rect 3164 272 3341 318
rect 3387 272 3564 318
rect 3610 272 3789 318
rect 3835 272 4014 318
rect 4060 272 4233 318
rect 4279 272 4290 318
rect 811 228 822 263
rect 2670 219 2728 272
rect 4446 219 4626 501
rect 4726 400 4737 446
rect 4783 400 4940 446
rect 4986 400 5144 446
rect 5190 400 5346 446
rect 5392 400 5553 446
rect 5599 400 5752 446
rect 5798 400 5959 446
rect 6005 400 6016 446
rect 4698 272 4709 318
rect 4755 272 4910 318
rect 4956 272 5134 318
rect 5180 272 5356 318
rect 5402 272 5584 318
rect 5630 272 5797 318
rect 5843 272 6019 318
rect 6065 272 6247 318
rect 6293 272 6304 318
rect 1202 187 1213 219
rect 262 82 273 128
rect 319 82 330 128
rect 843 173 1213 187
rect 1259 173 1661 219
rect 1707 173 2109 219
rect 2155 173 2557 219
rect 2603 173 2728 219
rect 2994 173 3005 219
rect 3051 173 3453 219
rect 3499 173 3901 219
rect 3947 173 4349 219
rect 4395 173 4797 219
rect 4843 173 5245 219
rect 5291 173 5693 219
rect 5739 173 6141 219
rect 6187 173 6198 219
rect 843 152 1270 173
rect 543 141 1270 152
rect 6365 141 6411 180
rect 543 123 888 141
rect 497 106 888 123
rect 262 60 330 82
rect 934 60 945 95
rect 0 49 945 60
rect 991 60 1002 95
rect 1426 81 1437 127
rect 1483 81 1494 127
rect 1426 60 1494 81
rect 1874 81 1885 127
rect 1931 81 1942 127
rect 1874 60 1942 81
rect 2322 81 2333 127
rect 2379 81 2390 127
rect 2322 60 2390 81
rect 2767 81 2781 127
rect 2827 81 2842 127
rect 2767 60 2842 81
rect 3218 81 3229 127
rect 3275 81 3286 127
rect 3218 60 3286 81
rect 3666 81 3677 127
rect 3723 81 3734 127
rect 3666 60 3734 81
rect 4114 81 4125 127
rect 4171 81 4182 127
rect 4114 60 4182 81
rect 4562 81 4573 127
rect 4619 81 4630 127
rect 4562 60 4630 81
rect 5010 81 5021 127
rect 5067 81 5078 127
rect 5010 60 5078 81
rect 5458 81 5469 127
rect 5515 81 5526 127
rect 5458 60 5526 81
rect 5906 81 5917 127
rect 5963 81 5974 127
rect 5906 60 5974 81
rect 6365 60 6411 95
rect 991 49 6496 60
rect 0 -60 6496 49
<< labels >>
flabel metal1 s 1138 354 2558 430 0 FreeSans 600 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 724 6496 844 0 FreeSans 600 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 6365 128 6411 180 0 FreeSans 600 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 5846 611 5914 676 0 FreeSans 600 0 0 0 Z
port 3 nsew default output
flabel metal1 s 74 354 318 430 0 FreeSans 600 0 0 0 EN
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 5438 611 5506 676 1 Z
port 3 nsew default output
rlabel metal1 s 5030 611 5098 676 1 Z
port 3 nsew default output
rlabel metal1 s 4626 611 4690 676 1 Z
port 3 nsew default output
rlabel metal1 s 4214 611 4282 676 1 Z
port 3 nsew default output
rlabel metal1 s 3806 611 3874 676 1 Z
port 3 nsew default output
rlabel metal1 s 3398 611 3466 676 1 Z
port 3 nsew default output
rlabel metal1 s 2990 611 3058 676 1 Z
port 3 nsew default output
rlabel metal1 s 2990 501 5914 611 1 Z
port 3 nsew default output
rlabel metal1 s 4446 219 4626 501 1 Z
port 3 nsew default output
rlabel metal1 s 2994 173 6198 219 1 Z
port 3 nsew default output
rlabel metal1 s 6061 657 6107 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5642 657 5710 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5234 657 5302 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4826 657 4894 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4418 657 4486 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4010 657 4078 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3602 657 3670 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3194 657 3262 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2786 657 2854 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2342 657 2410 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 657 1942 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 657 1534 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 657 1126 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 657 358 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6061 652 6107 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2786 652 2854 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2342 652 2410 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 652 1942 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 652 1534 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 652 1126 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6061 608 6107 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2786 608 2854 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2342 608 2410 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 608 1942 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 608 1534 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 608 1126 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6061 506 6107 608 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2786 506 2854 608 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6365 127 6411 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 127 330 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6365 95 6411 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5906 95 5974 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5458 95 5526 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5010 95 5078 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4562 95 4630 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4114 95 4182 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 95 3734 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 95 3286 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2767 95 2842 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 95 2390 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 95 1942 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 95 1494 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 95 330 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6365 60 6411 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5906 60 5974 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5458 60 5526 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5010 60 5078 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4562 60 4630 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4114 60 4182 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 60 3734 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 60 3286 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2767 60 2842 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 60 2390 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 60 1942 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 60 1494 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6496 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6496 784
string GDS_END 1440990
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1427948
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
