// Created Sat Aug 23 14:13:18 2025

module gf180mcu_fd_sc_mcu7t5v0__inv_1 (I, ZN, VDD, VNW, VPW, VSS);
  input  I;
  output ZN;
  inout  VDD;
  inout  VNW;
  inout  VPW;
  inout  VSS;
  // Functional behavior with power awareness
  assign ZN =  ~I;

  // Optional timing (edit tplh/tphl as needed)
endmodule

