magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 4100 1270
<< nmos >>
rect 190 210 250 380
rect 540 210 600 380
rect 710 210 770 380
rect 820 210 880 380
rect 1220 210 1280 380
rect 1430 210 1490 380
rect 1660 210 1720 380
rect 1770 210 1830 380
rect 1940 210 2000 380
rect 2050 210 2110 380
rect 2280 210 2340 380
rect 2490 210 2550 380
rect 2660 210 2720 380
rect 3040 210 3100 380
rect 3150 210 3210 380
rect 3320 210 3380 380
rect 3670 210 3730 380
rect 3840 210 3900 380
<< pmos >>
rect 190 720 250 1060
rect 510 720 570 1060
rect 680 720 740 1060
rect 850 720 910 1060
rect 1220 720 1280 1060
rect 1430 720 1490 1060
rect 1660 720 1720 1060
rect 1770 720 1830 1060
rect 1940 720 2000 1060
rect 2050 720 2110 1060
rect 2280 720 2340 1060
rect 2490 720 2550 1060
rect 2660 720 2720 1060
rect 3010 720 3070 1060
rect 3180 720 3240 1060
rect 3350 720 3410 1060
rect 3670 720 3730 1060
rect 3840 720 3900 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 440 278 540 380
rect 440 232 462 278
rect 508 232 540 278
rect 440 210 540 232
rect 600 303 710 380
rect 600 257 632 303
rect 678 257 710 303
rect 600 210 710 257
rect 770 210 820 380
rect 880 283 980 380
rect 880 237 912 283
rect 958 237 980 283
rect 880 210 980 237
rect 1120 283 1220 380
rect 1120 237 1142 283
rect 1188 237 1220 283
rect 1120 210 1220 237
rect 1280 210 1430 380
rect 1490 283 1660 380
rect 1490 237 1552 283
rect 1598 237 1660 283
rect 1490 210 1660 237
rect 1720 210 1770 380
rect 1830 278 1940 380
rect 1830 232 1862 278
rect 1908 232 1940 278
rect 1830 210 1940 232
rect 2000 210 2050 380
rect 2110 278 2280 380
rect 2110 232 2172 278
rect 2218 232 2280 278
rect 2110 210 2280 232
rect 2340 210 2490 380
rect 2550 303 2660 380
rect 2550 257 2582 303
rect 2628 257 2660 303
rect 2550 210 2660 257
rect 2720 318 2820 380
rect 2720 272 2752 318
rect 2798 272 2820 318
rect 2720 210 2820 272
rect 2940 318 3040 380
rect 2940 272 2962 318
rect 3008 272 3040 318
rect 2940 210 3040 272
rect 3100 210 3150 380
rect 3210 293 3320 380
rect 3210 247 3242 293
rect 3288 247 3320 293
rect 3210 210 3320 247
rect 3380 278 3480 380
rect 3380 232 3412 278
rect 3458 232 3480 278
rect 3380 210 3480 232
rect 3570 318 3670 380
rect 3570 272 3592 318
rect 3638 272 3670 318
rect 3570 210 3670 272
rect 3730 298 3840 380
rect 3730 252 3762 298
rect 3808 252 3840 298
rect 3730 210 3840 252
rect 3900 318 4000 380
rect 3900 272 3932 318
rect 3978 272 4000 318
rect 3900 210 4000 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 350 1060
rect 250 773 282 1007
rect 328 773 350 1007
rect 250 720 350 773
rect 410 1040 510 1060
rect 410 900 432 1040
rect 478 900 510 1040
rect 410 720 510 900
rect 570 1035 680 1060
rect 570 895 602 1035
rect 648 895 680 1035
rect 570 720 680 895
rect 740 1035 850 1060
rect 740 895 772 1035
rect 818 895 850 1035
rect 740 720 850 895
rect 910 1035 1010 1060
rect 910 895 942 1035
rect 988 895 1010 1035
rect 910 720 1010 895
rect 1120 1038 1220 1060
rect 1120 992 1142 1038
rect 1188 992 1220 1038
rect 1120 720 1220 992
rect 1280 720 1430 1060
rect 1490 1030 1660 1060
rect 1490 890 1552 1030
rect 1598 890 1660 1030
rect 1490 720 1660 890
rect 1720 720 1770 1060
rect 1830 1020 1940 1060
rect 1830 880 1862 1020
rect 1908 880 1940 1020
rect 1830 720 1940 880
rect 2000 720 2050 1060
rect 2110 1027 2280 1060
rect 2110 793 2172 1027
rect 2218 793 2280 1027
rect 2110 720 2280 793
rect 2340 720 2490 1060
rect 2550 1038 2660 1060
rect 2550 992 2582 1038
rect 2628 992 2660 1038
rect 2550 720 2660 992
rect 2720 1017 2820 1060
rect 2720 783 2752 1017
rect 2798 783 2820 1017
rect 2720 720 2820 783
rect 2910 1035 3010 1060
rect 2910 895 2932 1035
rect 2978 895 3010 1035
rect 2910 720 3010 895
rect 3070 1035 3180 1060
rect 3070 895 3102 1035
rect 3148 895 3180 1035
rect 3070 720 3180 895
rect 3240 1035 3350 1060
rect 3240 895 3272 1035
rect 3318 895 3350 1035
rect 3240 720 3350 895
rect 3410 1040 3510 1060
rect 3410 900 3442 1040
rect 3488 900 3510 1040
rect 3410 720 3510 900
rect 3570 1012 3670 1060
rect 3570 778 3592 1012
rect 3638 778 3670 1012
rect 3570 720 3670 778
rect 3730 1015 3840 1060
rect 3730 875 3762 1015
rect 3808 875 3840 1015
rect 3730 720 3840 875
rect 3900 1007 4000 1060
rect 3900 773 3932 1007
rect 3978 773 4000 1007
rect 3900 720 4000 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 462 232 508 278
rect 632 257 678 303
rect 912 237 958 283
rect 1142 237 1188 283
rect 1552 237 1598 283
rect 1862 232 1908 278
rect 2172 232 2218 278
rect 2582 257 2628 303
rect 2752 272 2798 318
rect 2962 272 3008 318
rect 3242 247 3288 293
rect 3412 232 3458 278
rect 3592 272 3638 318
rect 3762 252 3808 298
rect 3932 272 3978 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 432 900 478 1040
rect 602 895 648 1035
rect 772 895 818 1035
rect 942 895 988 1035
rect 1142 992 1188 1038
rect 1552 890 1598 1030
rect 1862 880 1908 1020
rect 2172 793 2218 1027
rect 2582 992 2628 1038
rect 2752 783 2798 1017
rect 2932 895 2978 1035
rect 3102 895 3148 1035
rect 3272 895 3318 1035
rect 3442 900 3488 1040
rect 3592 778 3638 1012
rect 3762 875 3808 1015
rect 3932 773 3978 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 550 118 700 140
rect 550 72 602 118
rect 648 72 700 118
rect 550 50 700 72
rect 790 118 940 140
rect 790 72 842 118
rect 888 72 940 118
rect 790 50 940 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
rect 2700 118 2850 140
rect 2700 72 2752 118
rect 2798 72 2850 118
rect 2700 50 2850 72
rect 2940 118 3090 140
rect 2940 72 2992 118
rect 3038 72 3090 118
rect 2940 50 3090 72
rect 3180 118 3330 140
rect 3180 72 3232 118
rect 3278 72 3330 118
rect 3180 50 3330 72
rect 3420 118 3570 140
rect 3420 72 3472 118
rect 3518 72 3570 118
rect 3420 50 3570 72
rect 3660 118 3810 140
rect 3660 72 3712 118
rect 3758 72 3810 118
rect 3660 50 3810 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 310 1198 460 1220
rect 310 1152 362 1198
rect 408 1152 460 1198
rect 310 1130 460 1152
rect 550 1198 700 1220
rect 550 1152 602 1198
rect 648 1152 700 1198
rect 550 1130 700 1152
rect 790 1198 940 1220
rect 790 1152 842 1198
rect 888 1152 940 1198
rect 790 1130 940 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
rect 1500 1198 1650 1220
rect 1500 1152 1552 1198
rect 1598 1152 1650 1198
rect 1500 1130 1650 1152
rect 1740 1198 1890 1220
rect 1740 1152 1792 1198
rect 1838 1152 1890 1198
rect 1740 1130 1890 1152
rect 1980 1198 2130 1220
rect 1980 1152 2032 1198
rect 2078 1152 2130 1198
rect 1980 1130 2130 1152
rect 2220 1198 2370 1220
rect 2220 1152 2272 1198
rect 2318 1152 2370 1198
rect 2220 1130 2370 1152
rect 2460 1198 2610 1220
rect 2460 1152 2512 1198
rect 2558 1152 2610 1198
rect 2460 1130 2610 1152
rect 2700 1198 2850 1220
rect 2700 1152 2752 1198
rect 2798 1152 2850 1198
rect 2700 1130 2850 1152
rect 2940 1198 3090 1220
rect 2940 1152 2992 1198
rect 3038 1152 3090 1198
rect 2940 1130 3090 1152
rect 3180 1198 3330 1220
rect 3180 1152 3232 1198
rect 3278 1152 3330 1198
rect 3180 1130 3330 1152
rect 3420 1198 3570 1220
rect 3420 1152 3472 1198
rect 3518 1152 3570 1198
rect 3420 1130 3570 1152
rect 3660 1198 3810 1220
rect 3660 1152 3712 1198
rect 3758 1152 3810 1198
rect 3660 1130 3810 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 602 72 648 118
rect 842 72 888 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
rect 2752 72 2798 118
rect 2992 72 3038 118
rect 3232 72 3278 118
rect 3472 72 3518 118
rect 3712 72 3758 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 362 1152 408 1198
rect 602 1152 648 1198
rect 842 1152 888 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
rect 1552 1152 1598 1198
rect 1792 1152 1838 1198
rect 2032 1152 2078 1198
rect 2272 1152 2318 1198
rect 2512 1152 2558 1198
rect 2752 1152 2798 1198
rect 2992 1152 3038 1198
rect 3232 1152 3278 1198
rect 3472 1152 3518 1198
rect 3712 1152 3758 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 510 1060 570 1110
rect 680 1060 740 1110
rect 850 1060 910 1110
rect 1220 1060 1280 1110
rect 1430 1060 1490 1110
rect 1660 1060 1720 1110
rect 1770 1060 1830 1110
rect 1940 1060 2000 1110
rect 2050 1060 2110 1110
rect 2280 1060 2340 1110
rect 2490 1060 2550 1110
rect 2660 1060 2720 1110
rect 3010 1060 3070 1110
rect 3180 1060 3240 1110
rect 3350 1060 3410 1110
rect 3670 1060 3730 1110
rect 3840 1060 3900 1110
rect 190 670 250 720
rect 140 643 250 670
rect 140 597 167 643
rect 213 597 250 643
rect 140 570 250 597
rect 190 380 250 570
rect 510 540 570 720
rect 680 700 740 720
rect 850 700 910 720
rect 680 673 800 700
rect 680 627 707 673
rect 753 627 800 673
rect 680 600 800 627
rect 850 673 990 700
rect 850 627 907 673
rect 953 627 990 673
rect 1220 670 1280 720
rect 1430 700 1490 720
rect 1360 673 1490 700
rect 850 600 990 627
rect 1200 643 1310 670
rect 510 513 630 540
rect 510 467 557 513
rect 603 467 630 513
rect 510 440 630 467
rect 680 450 740 600
rect 850 450 910 600
rect 1200 597 1237 643
rect 1283 597 1310 643
rect 1360 627 1387 673
rect 1433 670 1490 673
rect 1433 627 1460 670
rect 1360 600 1460 627
rect 1660 620 1720 720
rect 1770 700 1830 720
rect 1940 700 2000 720
rect 1770 630 2000 700
rect 2050 630 2110 720
rect 2280 700 2340 720
rect 2280 673 2400 700
rect 2280 670 2327 673
rect 1200 570 1310 597
rect 1510 570 1720 620
rect 540 380 600 440
rect 680 400 770 450
rect 710 380 770 400
rect 820 410 910 450
rect 820 380 880 410
rect 1220 380 1280 570
rect 1510 530 1570 570
rect 1390 503 1570 530
rect 1390 457 1427 503
rect 1473 457 1570 503
rect 1390 430 1570 457
rect 1620 498 1720 520
rect 1850 500 1910 630
rect 2050 580 2250 630
rect 2300 627 2327 670
rect 2373 627 2400 673
rect 2300 600 2400 627
rect 2490 590 2550 720
rect 2660 670 2720 720
rect 2660 643 2760 670
rect 2660 597 2687 643
rect 2733 597 2760 643
rect 2200 550 2250 580
rect 2470 563 2570 590
rect 1620 452 1647 498
rect 1693 452 1720 498
rect 1620 430 1720 452
rect 1430 380 1490 430
rect 1660 380 1720 430
rect 1770 480 1910 500
rect 2050 508 2150 530
rect 1770 473 2000 480
rect 1770 427 1807 473
rect 1853 427 2000 473
rect 1770 400 2000 427
rect 1770 380 1830 400
rect 1940 380 2000 400
rect 2050 462 2077 508
rect 2123 462 2150 508
rect 2200 523 2370 550
rect 2200 480 2287 523
rect 2050 440 2150 462
rect 2260 477 2287 480
rect 2333 477 2370 523
rect 2470 517 2497 563
rect 2543 517 2570 563
rect 2470 490 2570 517
rect 2660 570 2760 597
rect 2260 450 2370 477
rect 2050 380 2110 440
rect 2280 380 2340 450
rect 2490 380 2550 490
rect 2660 380 2720 570
rect 3010 510 3070 720
rect 2910 483 3070 510
rect 2910 437 2947 483
rect 2993 480 3070 483
rect 3180 670 3240 720
rect 3180 643 3280 670
rect 3180 597 3207 643
rect 3253 597 3280 643
rect 3180 570 3280 597
rect 2993 437 3100 480
rect 3180 450 3240 570
rect 3350 520 3410 720
rect 3670 610 3730 720
rect 3840 690 3900 720
rect 2910 410 3100 437
rect 3040 380 3100 410
rect 3150 400 3240 450
rect 3300 498 3410 520
rect 3620 583 3730 610
rect 3790 668 3900 690
rect 3790 622 3812 668
rect 3858 622 3900 668
rect 3790 600 3900 622
rect 3620 537 3647 583
rect 3693 537 3730 583
rect 3620 510 3730 537
rect 3300 452 3327 498
rect 3373 452 3410 498
rect 3300 430 3410 452
rect 3150 380 3210 400
rect 3320 380 3380 430
rect 3670 380 3730 510
rect 3840 380 3900 600
rect 190 160 250 210
rect 540 160 600 210
rect 710 160 770 210
rect 820 160 880 210
rect 1220 160 1280 210
rect 1430 160 1490 210
rect 1660 160 1720 210
rect 1770 160 1830 210
rect 1940 160 2000 210
rect 2050 160 2110 210
rect 2280 160 2340 210
rect 2490 160 2550 210
rect 2660 160 2720 210
rect 3040 160 3100 210
rect 3150 160 3210 210
rect 3320 160 3380 210
rect 3670 160 3730 210
rect 3840 160 3900 210
<< polycontact >>
rect 167 597 213 643
rect 707 627 753 673
rect 907 627 953 673
rect 557 467 603 513
rect 1237 597 1283 643
rect 1387 627 1433 673
rect 1427 457 1473 503
rect 2327 627 2373 673
rect 2687 597 2733 643
rect 1647 452 1693 498
rect 1807 427 1853 473
rect 2077 462 2123 508
rect 2287 477 2333 523
rect 2497 517 2543 563
rect 2947 437 2993 483
rect 3207 597 3253 643
rect 3812 622 3858 668
rect 3647 537 3693 583
rect 3327 452 3373 498
<< metal1 >>
rect 0 1198 4100 1270
rect 0 1152 112 1198
rect 158 1152 362 1198
rect 408 1152 602 1198
rect 648 1152 842 1198
rect 888 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1552 1198
rect 1598 1152 1792 1198
rect 1838 1152 2032 1198
rect 2078 1152 2272 1198
rect 2318 1152 2512 1198
rect 2558 1152 2752 1198
rect 2798 1152 2992 1198
rect 3038 1152 3232 1198
rect 3278 1152 3472 1198
rect 3518 1152 3712 1198
rect 3758 1152 4100 1198
rect 0 1130 4100 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 160 646 220 670
rect 160 594 164 646
rect 216 594 220 646
rect 160 570 220 594
rect 280 530 330 773
rect 430 1040 480 1060
rect 430 900 432 1040
rect 478 900 480 1040
rect 280 520 340 530
rect 280 516 360 520
rect 280 464 284 516
rect 336 464 360 516
rect 280 460 360 464
rect 280 400 340 460
rect 430 400 480 900
rect 600 1035 650 1060
rect 600 895 602 1035
rect 648 895 650 1035
rect 600 820 650 895
rect 770 1035 820 1130
rect 770 895 772 1035
rect 818 895 820 1035
rect 770 870 820 895
rect 940 1035 990 1060
rect 940 895 942 1035
rect 988 895 990 1035
rect 1140 1038 1190 1130
rect 1140 992 1142 1038
rect 1188 992 1190 1038
rect 1140 970 1190 992
rect 1520 1030 1630 1060
rect 1520 920 1552 1030
rect 940 820 990 895
rect 600 770 990 820
rect 1080 890 1552 920
rect 1598 890 1630 1030
rect 1080 860 1630 890
rect 1860 1020 1910 1130
rect 1860 880 1862 1020
rect 1908 880 1910 1020
rect 1080 680 1140 860
rect 1860 840 1910 880
rect 2140 1027 2250 1060
rect 2140 806 2172 1027
rect 2140 754 2164 806
rect 2218 793 2250 1027
rect 2580 1038 2630 1130
rect 2580 992 2582 1038
rect 2628 992 2630 1038
rect 2580 970 2630 992
rect 2750 1017 2800 1060
rect 2470 916 2570 920
rect 2470 864 2494 916
rect 2546 864 2570 916
rect 2470 860 2570 864
rect 2490 840 2550 860
rect 2216 754 2250 793
rect 2140 730 2250 754
rect 2750 783 2752 1017
rect 2798 790 2800 1017
rect 2930 1035 2980 1060
rect 2930 895 2932 1035
rect 2978 895 2980 1035
rect 2930 820 2980 895
rect 3100 1035 3150 1130
rect 3100 895 3102 1035
rect 3148 895 3150 1035
rect 3100 870 3150 895
rect 3270 1035 3320 1060
rect 3270 895 3272 1035
rect 3318 895 3320 1035
rect 3270 820 3320 895
rect 2798 783 2860 790
rect 2750 740 2860 783
rect 2930 770 3320 820
rect 3440 1040 3490 1060
rect 3440 900 3442 1040
rect 3488 900 3490 1040
rect 3440 840 3490 900
rect 3590 1012 3640 1060
rect 3440 790 3500 840
rect 680 676 780 680
rect 680 624 704 676
rect 756 624 780 676
rect 680 620 780 624
rect 880 676 1140 680
rect 880 624 904 676
rect 956 624 1140 676
rect 1360 673 2740 680
rect 880 620 1140 624
rect 1080 520 1140 620
rect 1210 646 1310 650
rect 1210 594 1234 646
rect 1286 594 1310 646
rect 1360 627 1387 673
rect 1433 627 2327 673
rect 2373 650 2740 673
rect 2373 646 2760 650
rect 2373 627 2684 646
rect 1360 620 2684 627
rect 1210 590 1310 594
rect 530 516 630 520
rect 530 464 554 516
rect 606 464 630 516
rect 530 460 630 464
rect 1080 460 1310 520
rect 1640 510 1700 620
rect 2070 510 2130 620
rect 2660 594 2684 620
rect 2736 594 2760 646
rect 2660 590 2760 594
rect 2470 566 2570 570
rect 2300 530 2360 560
rect 2260 526 2360 530
rect 2260 523 2304 526
rect 770 456 1030 460
rect 770 404 954 456
rect 1006 404 1030 456
rect 770 400 1030 404
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 400
rect 430 350 820 400
rect 280 272 282 318
rect 328 272 330 318
rect 630 340 820 350
rect 1250 350 1310 460
rect 1400 506 1500 510
rect 1400 454 1424 506
rect 1476 454 1500 506
rect 1400 450 1500 454
rect 1620 498 1720 510
rect 1620 452 1647 498
rect 1693 452 1720 498
rect 2050 508 2150 510
rect 1800 480 1860 490
rect 1620 450 1720 452
rect 1780 476 1880 480
rect 1780 424 1804 476
rect 1856 424 1880 476
rect 2050 462 2077 508
rect 2123 462 2150 508
rect 2260 477 2287 523
rect 2260 474 2304 477
rect 2356 474 2360 526
rect 2470 514 2494 566
rect 2546 514 2570 566
rect 2810 520 2860 740
rect 2910 646 3130 650
rect 2910 594 2934 646
rect 2986 594 3130 646
rect 2910 590 3130 594
rect 3180 646 3280 650
rect 3180 594 3204 646
rect 3256 594 3280 646
rect 3180 590 3280 594
rect 3450 590 3500 790
rect 3590 778 3592 1012
rect 3638 780 3640 1012
rect 3760 1015 3810 1130
rect 3760 875 3762 1015
rect 3808 875 3810 1015
rect 3930 1007 3980 1060
rect 3930 930 3932 1007
rect 3760 830 3810 875
rect 3920 906 3932 930
rect 3920 854 3924 906
rect 3920 830 3932 854
rect 3638 778 3880 780
rect 3590 776 3880 778
rect 3590 724 3804 776
rect 3856 724 3880 776
rect 3590 720 3880 724
rect 3930 773 3932 830
rect 3978 773 3980 1007
rect 3800 710 3860 720
rect 3810 668 3860 710
rect 3810 622 3812 668
rect 3858 622 3860 668
rect 2470 510 2570 514
rect 2260 470 2360 474
rect 2050 460 2150 462
rect 2300 460 2360 470
rect 2750 460 2860 520
rect 2920 486 3020 490
rect 1780 420 1880 424
rect 2300 410 2800 460
rect 2920 434 2944 486
rect 2996 434 3020 486
rect 2920 430 3020 434
rect 2140 386 2250 390
rect 630 303 680 340
rect 280 210 330 272
rect 460 278 510 300
rect 460 232 462 278
rect 508 232 510 278
rect 460 140 510 232
rect 630 257 632 303
rect 678 257 680 303
rect 630 210 680 257
rect 910 283 960 310
rect 910 237 912 283
rect 958 237 960 283
rect 910 140 960 237
rect 1140 283 1190 320
rect 1250 300 1630 350
rect 2140 334 2164 386
rect 2216 334 2250 386
rect 1140 237 1142 283
rect 1188 237 1190 283
rect 1140 140 1190 237
rect 1520 283 1630 300
rect 1520 237 1552 283
rect 1598 237 1630 283
rect 1520 210 1630 237
rect 1860 278 1910 300
rect 1860 232 1862 278
rect 1908 232 1910 278
rect 1860 140 1910 232
rect 2140 278 2250 334
rect 2140 232 2172 278
rect 2218 232 2250 278
rect 2140 210 2250 232
rect 2580 303 2630 360
rect 2580 257 2582 303
rect 2628 257 2630 303
rect 2580 140 2630 257
rect 2750 318 2800 410
rect 3070 400 3130 590
rect 3450 586 3720 590
rect 3450 534 3644 586
rect 3696 534 3720 586
rect 3450 530 3720 534
rect 3300 506 3400 510
rect 3300 454 3324 506
rect 3376 454 3400 506
rect 3300 452 3327 454
rect 3373 452 3400 454
rect 3300 450 3400 452
rect 3450 400 3500 530
rect 3810 440 3860 622
rect 2750 272 2752 318
rect 2798 272 2800 318
rect 2750 210 2800 272
rect 2960 318 3010 380
rect 3070 350 3500 400
rect 3590 390 3860 440
rect 2960 272 2962 318
rect 3008 272 3010 318
rect 2960 140 3010 272
rect 3240 293 3290 350
rect 3590 318 3640 390
rect 3240 247 3242 293
rect 3288 247 3290 293
rect 3240 210 3290 247
rect 3410 278 3460 300
rect 3410 232 3412 278
rect 3458 232 3460 278
rect 3410 140 3460 232
rect 3590 272 3592 318
rect 3638 272 3640 318
rect 3590 210 3640 272
rect 3760 298 3810 340
rect 3760 252 3762 298
rect 3808 252 3810 298
rect 3760 140 3810 252
rect 3930 318 3980 773
rect 3930 272 3932 318
rect 3978 272 3980 318
rect 3930 210 3980 272
rect 0 118 4100 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 602 118
rect 648 72 842 118
rect 888 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2752 118
rect 2798 72 2992 118
rect 3038 72 3232 118
rect 3278 72 3472 118
rect 3518 72 3712 118
rect 3758 72 4100 118
rect 0 0 4100 72
<< via1 >>
rect 164 643 216 646
rect 164 597 167 643
rect 167 597 213 643
rect 213 597 216 643
rect 164 594 216 597
rect 284 464 336 516
rect 2164 793 2172 806
rect 2172 793 2216 806
rect 2494 864 2546 916
rect 2164 754 2216 793
rect 704 673 756 676
rect 704 627 707 673
rect 707 627 753 673
rect 753 627 756 673
rect 704 624 756 627
rect 904 673 956 676
rect 904 627 907 673
rect 907 627 953 673
rect 953 627 956 673
rect 904 624 956 627
rect 1234 643 1286 646
rect 1234 597 1237 643
rect 1237 597 1283 643
rect 1283 597 1286 643
rect 1234 594 1286 597
rect 2684 643 2736 646
rect 554 513 606 516
rect 554 467 557 513
rect 557 467 603 513
rect 603 467 606 513
rect 554 464 606 467
rect 2684 597 2687 643
rect 2687 597 2733 643
rect 2733 597 2736 643
rect 2684 594 2736 597
rect 2304 523 2356 526
rect 954 404 1006 456
rect 1424 503 1476 506
rect 1424 457 1427 503
rect 1427 457 1473 503
rect 1473 457 1476 503
rect 1424 454 1476 457
rect 1804 473 1856 476
rect 1804 427 1807 473
rect 1807 427 1853 473
rect 1853 427 1856 473
rect 1804 424 1856 427
rect 2304 477 2333 523
rect 2333 477 2356 523
rect 2304 474 2356 477
rect 2494 563 2546 566
rect 2494 517 2497 563
rect 2497 517 2543 563
rect 2543 517 2546 563
rect 2494 514 2546 517
rect 2934 594 2986 646
rect 3204 643 3256 646
rect 3204 597 3207 643
rect 3207 597 3253 643
rect 3253 597 3256 643
rect 3204 594 3256 597
rect 3924 854 3932 906
rect 3932 854 3976 906
rect 3804 724 3856 776
rect 2944 483 2996 486
rect 2944 437 2947 483
rect 2947 437 2993 483
rect 2993 437 2996 483
rect 2944 434 2996 437
rect 2164 334 2216 386
rect 3644 583 3696 586
rect 3644 537 3647 583
rect 3647 537 3693 583
rect 3693 537 3696 583
rect 3644 534 3696 537
rect 3324 498 3376 506
rect 3324 454 3327 498
rect 3327 454 3373 498
rect 3373 454 3376 498
<< metal2 >>
rect 700 1010 3260 1070
rect 700 690 760 1010
rect 1420 890 2360 950
rect 2480 920 2560 930
rect 680 676 780 690
rect 150 650 230 660
rect 140 646 240 650
rect 140 594 164 646
rect 216 594 240 646
rect 680 624 704 676
rect 756 624 780 676
rect 680 610 780 624
rect 880 676 980 690
rect 880 624 904 676
rect 956 624 980 676
rect 1210 650 1310 660
rect 880 610 980 624
rect 1200 646 1320 650
rect 140 590 240 594
rect 1200 594 1234 646
rect 1286 594 1320 646
rect 1200 590 1320 594
rect 150 580 230 590
rect 1210 580 1310 590
rect 270 520 350 530
rect 530 520 630 530
rect 1420 520 1480 890
rect 2160 820 2220 830
rect 2150 806 2230 820
rect 2150 754 2164 806
rect 2216 754 2230 806
rect 2150 740 2230 754
rect 260 516 630 520
rect 260 464 284 516
rect 336 464 554 516
rect 606 464 630 516
rect 1410 510 1500 520
rect 1400 506 1500 510
rect 260 460 630 464
rect 270 450 350 460
rect 530 450 630 460
rect 930 460 1030 470
rect 930 456 1320 460
rect 550 260 610 450
rect 930 404 954 456
rect 1006 404 1320 456
rect 1400 454 1424 506
rect 1476 454 1500 506
rect 1800 490 1860 500
rect 1400 450 1500 454
rect 1410 440 1500 450
rect 1790 480 1870 490
rect 1790 476 1880 480
rect 930 400 1320 404
rect 930 390 1030 400
rect 1260 380 1320 400
rect 1790 424 1804 476
rect 1856 424 1880 476
rect 1790 420 1880 424
rect 1790 410 1870 420
rect 1790 380 1860 410
rect 2160 400 2220 740
rect 2300 540 2360 890
rect 2470 916 2900 920
rect 2470 864 2494 916
rect 2546 864 2900 916
rect 2470 860 2900 864
rect 2480 850 2560 860
rect 2490 580 2550 850
rect 2840 660 2900 860
rect 3200 660 3260 1010
rect 3910 910 3990 920
rect 3900 906 4000 910
rect 3900 854 3924 906
rect 3976 854 4000 906
rect 3900 850 4000 854
rect 3910 840 3990 850
rect 3790 780 3870 790
rect 3780 776 3880 780
rect 3780 724 3804 776
rect 3856 724 3880 776
rect 3780 720 3880 724
rect 3790 710 3870 720
rect 2670 650 2750 660
rect 2660 646 2760 650
rect 2660 594 2684 646
rect 2736 594 2760 646
rect 2660 590 2760 594
rect 2840 646 3010 660
rect 2840 594 2934 646
rect 2986 594 3010 646
rect 2840 590 3010 594
rect 2670 580 2750 590
rect 2910 580 3010 590
rect 3180 646 3280 660
rect 3180 594 3204 646
rect 3256 594 3280 646
rect 3180 580 3280 594
rect 3630 590 3710 600
rect 3600 586 3720 590
rect 2480 570 2560 580
rect 2470 566 2570 570
rect 2290 526 2370 540
rect 2290 474 2304 526
rect 2356 474 2370 526
rect 2470 514 2494 566
rect 2546 514 2570 566
rect 3600 534 3644 586
rect 3696 534 3720 586
rect 3600 530 3720 534
rect 3320 520 3380 530
rect 3630 520 3710 530
rect 2470 510 2570 514
rect 2480 500 2560 510
rect 3310 506 3390 520
rect 2290 460 2370 474
rect 2920 486 3020 500
rect 2300 450 2360 460
rect 2920 434 2944 486
rect 2996 434 3020 486
rect 2920 420 3020 434
rect 3310 454 3324 506
rect 3376 454 3390 506
rect 3310 430 3390 454
rect 2150 390 2230 400
rect 2920 390 3000 420
rect 1260 320 1860 380
rect 2140 386 3000 390
rect 2140 334 2164 386
rect 2216 334 3000 386
rect 2140 330 3000 334
rect 2150 320 2230 330
rect 3310 260 3370 430
rect 550 200 3370 260
<< labels >>
rlabel via1 s 1234 594 1286 646 4 D
port 1 nsew signal input
rlabel via1 s 3924 854 3976 906 4 Q
port 2 nsew signal output
rlabel via1 s 3804 724 3856 776 4 QN
port 3 nsew signal output
rlabel via1 s 3204 594 3256 646 4 SN
port 4 nsew signal output
rlabel via1 s 164 594 216 646 4 RN
port 5 nsew signal input
rlabel via1 s 2684 594 2736 646 4 CLK
port 6 nsew clock input
rlabel metal1 s 110 720 160 1270 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 770 870 820 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1140 970 1190 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1860 840 1910 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2580 970 2630 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3100 870 3150 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3760 830 3810 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 1130 4100 1270 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 460 0 510 300 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 910 0 960 310 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1140 0 1190 320 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1860 0 1910 300 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2580 0 2630 360 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2960 0 3010 380 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3410 0 3460 300 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3760 0 3810 340 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 0 4100 140 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal2 s 2670 580 2750 660 1 CLK
port 6 nsew clock input
rlabel metal2 s 2660 590 2760 650 1 CLK
port 6 nsew clock input
rlabel metal1 s 1640 450 1700 680 1 CLK
port 6 nsew clock input
rlabel metal1 s 1620 450 1720 510 1 CLK
port 6 nsew clock input
rlabel metal1 s 2070 460 2130 680 1 CLK
port 6 nsew clock input
rlabel metal1 s 2050 460 2150 510 1 CLK
port 6 nsew clock input
rlabel metal1 s 1360 620 2740 680 1 CLK
port 6 nsew clock input
rlabel metal1 s 2660 590 2760 650 1 CLK
port 6 nsew clock input
rlabel metal2 s 1210 580 1310 660 1 D
port 1 nsew signal input
rlabel metal2 s 1200 590 1320 650 1 D
port 1 nsew signal input
rlabel metal1 s 1210 590 1310 650 1 D
port 1 nsew signal input
rlabel metal2 s 3910 840 3990 920 1 Q
port 2 nsew signal output
rlabel metal2 s 3900 850 4000 910 1 Q
port 2 nsew signal output
rlabel metal1 s 3920 830 3980 930 1 Q
port 2 nsew signal output
rlabel metal1 s 3930 210 3980 1060 1 Q
port 2 nsew signal output
rlabel metal2 s 3790 710 3870 790 1 QN
port 3 nsew signal output
rlabel metal2 s 3780 720 3880 780 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 210 3640 440 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 720 3640 1060 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 390 3860 440 1 QN
port 3 nsew signal output
rlabel metal1 s 3810 390 3860 780 1 QN
port 3 nsew signal output
rlabel metal1 s 3800 710 3860 780 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 720 3880 780 1 QN
port 3 nsew signal output
rlabel metal2 s 150 580 230 660 1 RN
port 5 nsew signal input
rlabel metal2 s 140 590 240 650 1 RN
port 5 nsew signal input
rlabel metal1 s 160 570 220 670 1 RN
port 5 nsew signal input
rlabel via1 s 704 624 756 676 1 SN
port 4 nsew signal output
rlabel metal2 s 700 610 760 1070 1 SN
port 4 nsew signal output
rlabel metal2 s 680 610 780 690 1 SN
port 4 nsew signal output
rlabel metal2 s 3200 580 3260 1070 1 SN
port 4 nsew signal output
rlabel metal2 s 700 1010 3260 1070 1 SN
port 4 nsew signal output
rlabel metal2 s 3180 580 3280 660 1 SN
port 4 nsew signal output
rlabel metal1 s 680 620 780 680 1 SN
port 4 nsew signal output
rlabel metal1 s 3180 590 3280 650 1 SN
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 4100 1270
string GDS_END 252376
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 222302
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
