magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 4566 1094
<< pwell >>
rect -86 -86 4566 453
<< mvnmos >>
rect 124 156 244 272
rect 348 156 468 272
rect 516 156 636 272
rect 740 156 860 272
rect 908 156 1028 272
rect 1320 174 1440 332
rect 1632 174 1752 332
rect 2000 216 2120 332
rect 2224 216 2344 332
rect 2392 216 2512 332
rect 2692 216 2812 332
rect 2916 216 3036 332
rect 3140 216 3260 332
rect 3400 68 3520 332
rect 3624 68 3744 332
rect 4012 69 4132 333
rect 4236 69 4356 333
<< mvpmos >>
rect 144 652 244 852
rect 368 652 468 852
rect 526 652 626 852
rect 750 652 850 852
rect 918 652 1018 852
rect 1448 573 1548 849
rect 1652 573 1752 849
rect 2166 652 2266 852
rect 2370 652 2470 852
rect 2518 652 2618 852
rect 2722 652 2822 852
rect 2926 652 3026 852
rect 3140 652 3240 852
rect 3400 573 3500 939
rect 3604 573 3704 939
rect 4022 574 4122 940
rect 4233 574 4333 940
<< mvndiff >>
rect 1232 319 1320 332
rect 1232 273 1245 319
rect 1291 273 1320 319
rect 36 215 124 272
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 272
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 272
rect 636 215 740 272
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 272
rect 1028 156 1160 272
rect 1232 174 1320 273
rect 1440 174 1632 332
rect 1752 319 1840 332
rect 1752 273 1781 319
rect 1827 273 1840 319
rect 1752 174 1840 273
rect 1912 275 2000 332
rect 1912 229 1925 275
rect 1971 229 2000 275
rect 1912 216 2000 229
rect 2120 319 2224 332
rect 2120 273 2149 319
rect 2195 273 2224 319
rect 2120 216 2224 273
rect 2344 216 2392 332
rect 2512 216 2692 332
rect 2812 319 2916 332
rect 2812 273 2841 319
rect 2887 273 2916 319
rect 2812 216 2916 273
rect 3036 319 3140 332
rect 3036 273 3065 319
rect 3111 273 3140 319
rect 3036 216 3140 273
rect 3260 216 3400 332
rect 1088 113 1160 156
rect 1088 67 1101 113
rect 1147 67 1160 113
rect 1088 54 1160 67
rect 1500 113 1572 174
rect 1500 67 1513 113
rect 1559 67 1572 113
rect 1500 54 1572 67
rect 2572 126 2632 216
rect 2561 118 2632 126
rect 2561 113 2633 118
rect 2561 67 2574 113
rect 2620 67 2633 113
rect 3320 68 3400 216
rect 3520 307 3624 332
rect 3520 167 3549 307
rect 3595 167 3624 307
rect 3520 68 3624 167
rect 3744 309 3832 332
rect 3744 169 3773 309
rect 3819 169 3832 309
rect 3744 68 3832 169
rect 3924 309 4012 333
rect 3924 169 3937 309
rect 3983 169 4012 309
rect 3924 69 4012 169
rect 4132 320 4236 333
rect 4132 180 4161 320
rect 4207 180 4236 320
rect 4132 69 4236 180
rect 4356 222 4444 333
rect 4356 82 4385 222
rect 4431 82 4444 222
rect 4356 69 4444 82
rect 2561 54 2633 67
<< mvpdiff >>
rect 56 839 144 852
rect 56 699 69 839
rect 115 699 144 839
rect 56 652 144 699
rect 244 839 368 852
rect 244 699 273 839
rect 319 699 368 839
rect 244 652 368 699
rect 468 652 526 852
rect 626 839 750 852
rect 626 699 675 839
rect 721 699 750 839
rect 626 652 750 699
rect 850 652 918 852
rect 1018 838 1106 852
rect 3320 852 3400 939
rect 1018 792 1047 838
rect 1093 792 1106 838
rect 1018 652 1106 792
rect 1360 632 1448 849
rect 1360 586 1373 632
rect 1419 586 1448 632
rect 1360 573 1448 586
rect 1548 827 1652 849
rect 1548 781 1577 827
rect 1623 781 1652 827
rect 1548 573 1652 781
rect 1752 632 1840 849
rect 2078 746 2166 852
rect 2078 700 2091 746
rect 2137 700 2166 746
rect 2078 652 2166 700
rect 2266 839 2370 852
rect 2266 699 2295 839
rect 2341 699 2370 839
rect 2266 652 2370 699
rect 2470 652 2518 852
rect 2618 839 2722 852
rect 2618 699 2647 839
rect 2693 699 2722 839
rect 2618 652 2722 699
rect 2822 839 2926 852
rect 2822 699 2851 839
rect 2897 699 2926 839
rect 2822 652 2926 699
rect 3026 839 3140 852
rect 3026 699 3065 839
rect 3111 699 3140 839
rect 3026 652 3140 699
rect 3240 652 3400 852
rect 1752 586 1781 632
rect 1827 586 1840 632
rect 1752 573 1840 586
rect 3320 573 3400 652
rect 3500 871 3604 939
rect 3500 731 3529 871
rect 3575 731 3604 871
rect 3500 573 3604 731
rect 3704 839 3792 939
rect 3704 699 3733 839
rect 3779 699 3792 839
rect 3704 573 3792 699
rect 3934 927 4022 940
rect 3934 787 3947 927
rect 3993 787 4022 927
rect 3934 574 4022 787
rect 4122 839 4233 940
rect 4122 699 4158 839
rect 4204 699 4233 839
rect 4122 574 4233 699
rect 4333 927 4421 940
rect 4333 787 4362 927
rect 4408 787 4421 927
rect 4333 574 4421 787
<< mvndiffc >>
rect 1245 273 1291 319
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1781 273 1827 319
rect 1925 229 1971 275
rect 2149 273 2195 319
rect 2841 273 2887 319
rect 3065 273 3111 319
rect 1101 67 1147 113
rect 1513 67 1559 113
rect 2574 67 2620 113
rect 3549 167 3595 307
rect 3773 169 3819 309
rect 3937 169 3983 309
rect 4161 180 4207 320
rect 4385 82 4431 222
<< mvpdiffc >>
rect 69 699 115 839
rect 273 699 319 839
rect 675 699 721 839
rect 1047 792 1093 838
rect 1373 586 1419 632
rect 1577 781 1623 827
rect 2091 700 2137 746
rect 2295 699 2341 839
rect 2647 699 2693 839
rect 2851 699 2897 839
rect 3065 699 3111 839
rect 1781 586 1827 632
rect 3529 731 3575 871
rect 3733 699 3779 839
rect 3947 787 3993 927
rect 4158 699 4204 839
rect 4362 787 4408 927
<< polysilicon >>
rect 144 944 850 984
rect 144 852 244 944
rect 368 852 468 896
rect 526 852 626 896
rect 750 852 850 944
rect 1652 944 3026 984
rect 918 852 1018 896
rect 1448 849 1548 893
rect 1652 849 1752 944
rect 2166 852 2266 896
rect 2370 852 2470 944
rect 2518 852 2618 896
rect 2722 852 2822 896
rect 2926 852 3026 944
rect 3400 939 3500 983
rect 3604 939 3704 983
rect 4022 940 4122 984
rect 4233 940 4333 984
rect 3140 852 3240 896
rect 144 502 244 652
rect 144 456 157 502
rect 203 456 244 502
rect 144 316 244 456
rect 368 502 468 652
rect 526 513 626 652
rect 750 608 850 652
rect 918 515 1018 652
rect 368 456 381 502
rect 427 456 468 502
rect 368 316 468 456
rect 520 502 626 513
rect 520 456 533 502
rect 579 456 626 502
rect 520 436 626 456
rect 908 502 1018 515
rect 908 456 921 502
rect 967 456 1018 502
rect 520 364 860 436
rect 124 272 244 316
rect 348 272 468 316
rect 516 272 636 316
rect 740 272 860 364
rect 908 316 1018 456
rect 1448 502 1548 573
rect 1448 456 1486 502
rect 1532 456 1548 502
rect 1448 432 1548 456
rect 1320 392 1548 432
rect 1652 502 1752 573
rect 1652 456 1665 502
rect 1711 456 1752 502
rect 1320 332 1440 392
rect 1652 376 1752 456
rect 2166 502 2266 652
rect 2370 608 2470 652
rect 2166 456 2179 502
rect 2225 456 2266 502
rect 2518 502 2618 652
rect 2722 608 2822 652
rect 2722 515 2812 608
rect 2518 464 2559 502
rect 2166 451 2266 456
rect 2392 456 2559 464
rect 2605 456 2618 502
rect 2166 392 2344 451
rect 1632 332 1752 376
rect 2000 332 2120 376
rect 2224 332 2344 392
rect 2392 392 2618 456
rect 2692 502 2812 515
rect 2692 456 2705 502
rect 2751 456 2812 502
rect 2392 332 2512 392
rect 2692 332 2812 456
rect 2926 464 3026 652
rect 3140 571 3240 652
rect 3140 525 3157 571
rect 3203 525 3240 571
rect 3140 512 3240 525
rect 3400 502 3500 573
rect 2926 424 3260 464
rect 2916 332 3036 376
rect 3140 332 3260 424
rect 3400 456 3441 502
rect 3487 456 3500 502
rect 3400 376 3500 456
rect 3604 502 3704 573
rect 3604 456 3617 502
rect 3663 456 3704 502
rect 3604 443 3704 456
rect 3624 376 3704 443
rect 3823 502 3923 515
rect 3823 456 3836 502
rect 3882 496 3923 502
rect 4022 496 4122 574
rect 4233 496 4333 574
rect 3882 456 4333 496
rect 3823 424 4333 456
rect 3400 332 3520 376
rect 3624 332 3744 376
rect 4012 333 4132 424
rect 4236 377 4333 424
rect 4236 333 4356 377
rect 908 272 1028 316
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1320 130 1440 174
rect 124 24 636 64
rect 1632 96 1752 174
rect 2000 96 2120 216
rect 2224 183 2344 216
rect 2224 137 2285 183
rect 2331 137 2344 183
rect 2392 172 2512 216
rect 2224 124 2344 137
rect 2692 172 2812 216
rect 2916 183 3036 216
rect 1632 24 2120 96
rect 2916 137 2957 183
rect 3003 137 3036 183
rect 3140 172 3260 216
rect 2916 124 3036 137
rect 3400 24 3520 68
rect 3624 24 3744 68
rect 4012 25 4132 69
rect 4236 25 4356 69
<< polycontact >>
rect 157 456 203 502
rect 381 456 427 502
rect 533 456 579 502
rect 921 456 967 502
rect 1486 456 1532 502
rect 1665 456 1711 502
rect 2179 456 2225 502
rect 2559 456 2605 502
rect 2705 456 2751 502
rect 3157 525 3203 571
rect 3441 456 3487 502
rect 3617 456 3663 502
rect 3836 456 3882 502
rect 2285 137 2331 183
rect 2957 137 3003 183
<< metal1 >>
rect 0 927 4480 1098
rect 0 918 3947 927
rect 69 839 115 850
rect 69 642 115 699
rect 273 839 319 918
rect 273 688 319 699
rect 675 839 1001 850
rect 721 804 1001 839
rect 675 688 721 699
rect 955 735 1001 804
rect 1047 838 1093 918
rect 1047 781 1093 792
rect 1566 827 1634 918
rect 1566 781 1577 827
rect 1623 781 1634 827
rect 2295 839 2341 850
rect 2091 746 2137 757
rect 955 700 2091 735
rect 955 689 2137 700
rect 69 596 579 642
rect 30 502 203 542
rect 30 456 157 502
rect 30 445 203 456
rect 366 502 427 542
rect 366 456 381 502
rect 30 354 82 445
rect 366 354 427 456
rect 533 502 579 596
rect 1373 632 1711 643
rect 1419 597 1711 632
rect 1373 575 1419 586
rect 533 308 579 456
rect 814 502 967 542
rect 814 456 921 502
rect 814 445 967 456
rect 1486 502 1538 542
rect 1532 456 1538 502
rect 814 354 866 445
rect 1486 354 1538 456
rect 1665 502 1711 597
rect 49 262 579 308
rect 1245 319 1291 330
rect 1665 308 1711 456
rect 1291 273 1711 308
rect 1245 262 1711 273
rect 1781 632 1827 643
rect 1781 513 1827 586
rect 1781 502 2225 513
rect 1781 456 2179 502
rect 1781 445 2225 456
rect 1781 319 1827 445
rect 2295 399 2341 699
rect 2647 839 2693 918
rect 3529 871 3575 918
rect 2647 688 2693 699
rect 2851 839 2897 850
rect 2851 605 2897 699
rect 2559 559 2897 605
rect 2559 502 2605 559
rect 2559 445 2605 456
rect 2705 502 2751 513
rect 2705 399 2751 456
rect 2295 353 2751 399
rect 2295 330 2341 353
rect 2149 319 2341 330
rect 1781 262 1827 273
rect 1925 275 1971 286
rect 49 215 95 262
rect 2195 273 2341 319
rect 2149 262 2341 273
rect 2841 319 2897 559
rect 2887 273 2897 319
rect 2841 262 2897 273
rect 3065 839 3111 850
rect 3529 720 3575 731
rect 3733 839 3779 850
rect 3065 674 3111 699
rect 3993 918 4362 927
rect 3947 776 3993 787
rect 4158 839 4226 850
rect 3065 628 3579 674
rect 3065 319 3111 628
rect 3065 262 3111 273
rect 3157 571 3203 582
rect 665 216 711 226
rect 1925 216 1971 229
rect 3157 216 3203 525
rect 3441 502 3487 513
rect 3533 502 3579 628
rect 3733 513 3779 699
rect 4204 699 4226 839
rect 4408 918 4480 927
rect 4362 776 4408 787
rect 3733 502 3882 513
rect 3533 456 3617 502
rect 3663 456 3674 502
rect 3733 456 3836 502
rect 3441 410 3487 456
rect 3733 445 3882 456
rect 3733 410 3819 445
rect 3441 364 3819 410
rect 665 215 1971 216
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 711 170 1971 215
rect 2274 183 3203 216
rect 665 158 711 169
rect 2274 137 2285 183
rect 2331 170 2957 183
rect 2331 137 2342 170
rect 2946 137 2957 170
rect 3003 137 3203 183
rect 3549 307 3595 318
rect 1101 113 1147 124
rect 0 67 1101 90
rect 1513 113 1559 124
rect 1147 67 1513 90
rect 2574 113 2620 124
rect 1559 67 2574 90
rect 3549 90 3595 167
rect 3773 309 3819 364
rect 4158 320 4226 699
rect 3773 158 3819 169
rect 3937 309 3983 320
rect 4158 180 4161 320
rect 4207 180 4226 320
rect 4158 169 4226 180
rect 4385 222 4431 233
rect 3937 90 3983 169
rect 2620 82 4385 90
rect 4431 82 4480 90
rect 2620 67 4480 82
rect 0 -90 4480 67
<< labels >>
flabel metal1 s 1486 354 1538 542 0 FreeSans 200 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 814 445 967 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4158 169 4226 850 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 30 445 203 542 0 FreeSans 200 0 0 0 SE
port 2 nsew default input
flabel metal1 s 366 354 427 542 0 FreeSans 200 0 0 0 SI
port 3 nsew default input
flabel metal1 s 0 918 4480 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3937 318 3983 320 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 814 354 866 445 1 D
port 1 nsew default input
rlabel metal1 s 30 354 82 445 1 SE
port 2 nsew default input
rlabel metal1 s 4362 781 4408 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 781 3993 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 781 3575 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2647 781 2693 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1566 781 1634 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1047 781 1093 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 781 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4362 776 4408 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 776 3993 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 776 3575 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2647 776 2693 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 776 319 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 720 3575 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2647 720 2693 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 720 319 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2647 688 2693 720 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 688 319 720 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3937 233 3983 318 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 233 3595 318 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4385 215 4431 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 215 3983 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 215 3595 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4385 124 4431 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 124 3983 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 124 3595 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 124 330 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4385 90 4431 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 90 3983 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 90 3595 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2574 90 2620 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1513 90 1559 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1101 90 1147 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 124 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4480 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4480 1008
string GDS_END 322628
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 312722
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
