magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 85 29129 22775 29790
rect 85 29053 23905 29129
rect 1342 27025 23905 29053
rect 1342 25454 23709 27025
rect 1342 23867 23707 25454
rect 1216 17407 22310 19961
rect 22338 18379 23707 19961
rect 22338 17923 23923 18379
rect 22338 17407 23905 17923
rect 22338 17406 22926 17407
rect 22827 14326 23842 15917
rect 22992 9181 23846 10665
rect 22880 8391 23846 9181
rect 22992 8114 23846 8391
rect 22861 7037 23846 7493
<< pwell >>
rect 239 89663 23775 89695
rect 239 30119 23775 30151
<< mvnmos >>
rect 23332 22316 23452 23678
rect 23332 20312 23452 21674
rect 23292 17142 23412 17256
rect 23516 17142 23636 17256
rect 23243 13889 23363 14165
rect 23467 13889 23587 14165
rect 23247 10804 23367 12504
rect 23471 10804 23591 12504
<< mvpmos >>
rect 361 29194 834 29649
rect 980 29194 1453 29649
rect 1599 29194 2072 29649
rect 2218 29194 2691 29649
rect 2837 29194 3310 29649
rect 3456 29194 3929 29649
rect 4075 29194 4548 29649
rect 4694 29194 5167 29649
rect 5313 29194 5786 29649
rect 5932 29194 6405 29649
rect 6551 29194 7024 29649
rect 7170 29194 7643 29649
rect 7789 29194 8262 29649
rect 8408 29194 8881 29649
rect 9027 29194 9500 29649
rect 9646 29194 10119 29649
rect 10265 29194 10738 29649
rect 10884 29194 11357 29649
rect 11503 29194 11976 29649
rect 12122 29194 12595 29649
rect 12741 29194 13214 29649
rect 13360 29194 13833 29649
rect 13979 29194 14452 29649
rect 14598 29194 15071 29649
rect 15217 29194 15690 29649
rect 15836 29194 16309 29649
rect 16455 29194 16928 29649
rect 17074 29194 17547 29649
rect 17693 29194 18166 29649
rect 18312 29194 18785 29649
rect 18931 29194 19404 29649
rect 19550 29194 20023 29649
rect 20169 29194 20642 29649
rect 20788 29194 21261 29649
rect 21407 29194 21880 29649
rect 22026 29194 22499 29649
rect 23220 27950 23340 28632
rect 23444 27950 23564 28632
rect 23220 27175 23340 27857
rect 23444 27175 23564 27857
rect 23334 25594 23454 26956
rect 23332 24007 23452 25369
rect 23332 18457 23452 19819
rect 23263 17547 23383 17844
rect 23515 17547 23635 17844
rect 23243 14469 23363 15171
rect 23467 14469 23587 15171
rect 23247 8395 23367 10523
rect 23471 8395 23591 10523
<< mvndiff >>
rect 23244 23665 23332 23678
rect 23244 23619 23257 23665
rect 23303 23619 23332 23665
rect 23244 23557 23332 23619
rect 23244 23511 23257 23557
rect 23303 23511 23332 23557
rect 23244 23449 23332 23511
rect 23244 23403 23257 23449
rect 23303 23403 23332 23449
rect 23244 23341 23332 23403
rect 23244 23295 23257 23341
rect 23303 23295 23332 23341
rect 23244 23233 23332 23295
rect 23244 23187 23257 23233
rect 23303 23187 23332 23233
rect 23244 23125 23332 23187
rect 23244 23079 23257 23125
rect 23303 23079 23332 23125
rect 23244 23017 23332 23079
rect 23244 22971 23257 23017
rect 23303 22971 23332 23017
rect 23244 22910 23332 22971
rect 23244 22864 23257 22910
rect 23303 22864 23332 22910
rect 23244 22803 23332 22864
rect 23244 22757 23257 22803
rect 23303 22757 23332 22803
rect 23244 22696 23332 22757
rect 23244 22650 23257 22696
rect 23303 22650 23332 22696
rect 23244 22589 23332 22650
rect 23244 22543 23257 22589
rect 23303 22543 23332 22589
rect 23244 22482 23332 22543
rect 23244 22436 23257 22482
rect 23303 22436 23332 22482
rect 23244 22375 23332 22436
rect 23244 22329 23257 22375
rect 23303 22329 23332 22375
rect 23244 22316 23332 22329
rect 23452 23665 23540 23678
rect 23452 23619 23481 23665
rect 23527 23619 23540 23665
rect 23452 23557 23540 23619
rect 23452 23511 23481 23557
rect 23527 23511 23540 23557
rect 23452 23449 23540 23511
rect 23452 23403 23481 23449
rect 23527 23403 23540 23449
rect 23452 23341 23540 23403
rect 23452 23295 23481 23341
rect 23527 23295 23540 23341
rect 23452 23233 23540 23295
rect 23452 23187 23481 23233
rect 23527 23187 23540 23233
rect 23452 23125 23540 23187
rect 23452 23079 23481 23125
rect 23527 23079 23540 23125
rect 23452 23017 23540 23079
rect 23452 22971 23481 23017
rect 23527 22971 23540 23017
rect 23452 22910 23540 22971
rect 23452 22864 23481 22910
rect 23527 22864 23540 22910
rect 23452 22803 23540 22864
rect 23452 22757 23481 22803
rect 23527 22757 23540 22803
rect 23452 22696 23540 22757
rect 23452 22650 23481 22696
rect 23527 22650 23540 22696
rect 23452 22589 23540 22650
rect 23452 22543 23481 22589
rect 23527 22543 23540 22589
rect 23452 22482 23540 22543
rect 23452 22436 23481 22482
rect 23527 22436 23540 22482
rect 23452 22375 23540 22436
rect 23452 22329 23481 22375
rect 23527 22329 23540 22375
rect 23452 22316 23540 22329
rect 23244 21661 23332 21674
rect 23244 21615 23257 21661
rect 23303 21615 23332 21661
rect 23244 21553 23332 21615
rect 23244 21507 23257 21553
rect 23303 21507 23332 21553
rect 23244 21445 23332 21507
rect 23244 21399 23257 21445
rect 23303 21399 23332 21445
rect 23244 21337 23332 21399
rect 23244 21291 23257 21337
rect 23303 21291 23332 21337
rect 23244 21229 23332 21291
rect 23244 21183 23257 21229
rect 23303 21183 23332 21229
rect 23244 21121 23332 21183
rect 23244 21075 23257 21121
rect 23303 21075 23332 21121
rect 23244 21013 23332 21075
rect 23244 20967 23257 21013
rect 23303 20967 23332 21013
rect 23244 20906 23332 20967
rect 23244 20860 23257 20906
rect 23303 20860 23332 20906
rect 23244 20799 23332 20860
rect 23244 20753 23257 20799
rect 23303 20753 23332 20799
rect 23244 20692 23332 20753
rect 23244 20646 23257 20692
rect 23303 20646 23332 20692
rect 23244 20585 23332 20646
rect 23244 20539 23257 20585
rect 23303 20539 23332 20585
rect 23244 20478 23332 20539
rect 23244 20432 23257 20478
rect 23303 20432 23332 20478
rect 23244 20371 23332 20432
rect 23244 20325 23257 20371
rect 23303 20325 23332 20371
rect 23244 20312 23332 20325
rect 23452 21661 23540 21674
rect 23452 21615 23481 21661
rect 23527 21615 23540 21661
rect 23452 21553 23540 21615
rect 23452 21507 23481 21553
rect 23527 21507 23540 21553
rect 23452 21445 23540 21507
rect 23452 21399 23481 21445
rect 23527 21399 23540 21445
rect 23452 21337 23540 21399
rect 23452 21291 23481 21337
rect 23527 21291 23540 21337
rect 23452 21229 23540 21291
rect 23452 21183 23481 21229
rect 23527 21183 23540 21229
rect 23452 21121 23540 21183
rect 23452 21075 23481 21121
rect 23527 21075 23540 21121
rect 23452 21013 23540 21075
rect 23452 20967 23481 21013
rect 23527 20967 23540 21013
rect 23452 20906 23540 20967
rect 23452 20860 23481 20906
rect 23527 20860 23540 20906
rect 23452 20799 23540 20860
rect 23452 20753 23481 20799
rect 23527 20753 23540 20799
rect 23452 20692 23540 20753
rect 23452 20646 23481 20692
rect 23527 20646 23540 20692
rect 23452 20585 23540 20646
rect 23452 20539 23481 20585
rect 23527 20539 23540 20585
rect 23452 20478 23540 20539
rect 23452 20432 23481 20478
rect 23527 20432 23540 20478
rect 23452 20371 23540 20432
rect 23452 20325 23481 20371
rect 23527 20325 23540 20371
rect 23452 20312 23540 20325
rect 23204 17222 23292 17256
rect 23204 17176 23217 17222
rect 23263 17176 23292 17222
rect 23204 17142 23292 17176
rect 23412 17222 23516 17256
rect 23412 17176 23441 17222
rect 23487 17176 23516 17222
rect 23412 17142 23516 17176
rect 23636 17222 23724 17256
rect 23636 17176 23665 17222
rect 23711 17176 23724 17222
rect 23636 17142 23724 17176
rect 23155 14152 23243 14165
rect 23155 13902 23168 14152
rect 23214 13902 23243 14152
rect 23155 13889 23243 13902
rect 23363 14152 23467 14165
rect 23363 13902 23392 14152
rect 23438 13902 23467 14152
rect 23363 13889 23467 13902
rect 23587 14152 23675 14165
rect 23587 13902 23616 14152
rect 23662 13902 23675 14152
rect 23587 13889 23675 13902
rect 23159 12491 23247 12504
rect 23159 10817 23172 12491
rect 23218 10817 23247 12491
rect 23159 10804 23247 10817
rect 23367 12491 23471 12504
rect 23367 10817 23396 12491
rect 23442 10817 23471 12491
rect 23367 10804 23471 10817
rect 23591 12491 23679 12504
rect 23591 10817 23620 12491
rect 23666 10817 23679 12491
rect 23591 10804 23679 10817
<< mvpdiff >>
rect 221 29604 361 29649
rect 221 29558 265 29604
rect 311 29558 361 29604
rect 221 29286 361 29558
rect 221 29240 265 29286
rect 311 29240 361 29286
rect 221 29194 361 29240
rect 834 29604 980 29649
rect 834 29558 884 29604
rect 930 29558 980 29604
rect 834 29286 980 29558
rect 834 29240 884 29286
rect 930 29240 980 29286
rect 834 29194 980 29240
rect 1453 29604 1599 29649
rect 1453 29558 1503 29604
rect 1549 29558 1599 29604
rect 1453 29286 1599 29558
rect 1453 29240 1503 29286
rect 1549 29240 1599 29286
rect 1453 29194 1599 29240
rect 2072 29604 2218 29649
rect 2072 29558 2122 29604
rect 2168 29558 2218 29604
rect 2072 29286 2218 29558
rect 2072 29240 2122 29286
rect 2168 29240 2218 29286
rect 2072 29194 2218 29240
rect 2691 29604 2837 29649
rect 2691 29558 2741 29604
rect 2787 29558 2837 29604
rect 2691 29286 2837 29558
rect 2691 29240 2741 29286
rect 2787 29240 2837 29286
rect 2691 29194 2837 29240
rect 3310 29604 3456 29649
rect 3310 29558 3360 29604
rect 3406 29558 3456 29604
rect 3310 29286 3456 29558
rect 3310 29240 3360 29286
rect 3406 29240 3456 29286
rect 3310 29194 3456 29240
rect 3929 29604 4075 29649
rect 3929 29558 3979 29604
rect 4025 29558 4075 29604
rect 3929 29286 4075 29558
rect 3929 29240 3979 29286
rect 4025 29240 4075 29286
rect 3929 29194 4075 29240
rect 4548 29604 4694 29649
rect 4548 29558 4598 29604
rect 4644 29558 4694 29604
rect 4548 29286 4694 29558
rect 4548 29240 4598 29286
rect 4644 29240 4694 29286
rect 4548 29194 4694 29240
rect 5167 29604 5313 29649
rect 5167 29558 5217 29604
rect 5263 29558 5313 29604
rect 5167 29286 5313 29558
rect 5167 29240 5217 29286
rect 5263 29240 5313 29286
rect 5167 29194 5313 29240
rect 5786 29604 5932 29649
rect 5786 29558 5836 29604
rect 5882 29558 5932 29604
rect 5786 29286 5932 29558
rect 5786 29240 5836 29286
rect 5882 29240 5932 29286
rect 5786 29194 5932 29240
rect 6405 29604 6551 29649
rect 6405 29558 6455 29604
rect 6501 29558 6551 29604
rect 6405 29286 6551 29558
rect 6405 29240 6455 29286
rect 6501 29240 6551 29286
rect 6405 29194 6551 29240
rect 7024 29604 7170 29649
rect 7024 29558 7074 29604
rect 7120 29558 7170 29604
rect 7024 29286 7170 29558
rect 7024 29240 7074 29286
rect 7120 29240 7170 29286
rect 7024 29194 7170 29240
rect 7643 29604 7789 29649
rect 7643 29558 7693 29604
rect 7739 29558 7789 29604
rect 7643 29286 7789 29558
rect 7643 29240 7693 29286
rect 7739 29240 7789 29286
rect 7643 29194 7789 29240
rect 8262 29604 8408 29649
rect 8262 29558 8312 29604
rect 8358 29558 8408 29604
rect 8262 29286 8408 29558
rect 8262 29240 8312 29286
rect 8358 29240 8408 29286
rect 8262 29194 8408 29240
rect 8881 29604 9027 29649
rect 8881 29558 8931 29604
rect 8977 29558 9027 29604
rect 8881 29286 9027 29558
rect 8881 29240 8931 29286
rect 8977 29240 9027 29286
rect 8881 29194 9027 29240
rect 9500 29604 9646 29649
rect 9500 29558 9550 29604
rect 9596 29558 9646 29604
rect 9500 29286 9646 29558
rect 9500 29240 9550 29286
rect 9596 29240 9646 29286
rect 9500 29194 9646 29240
rect 10119 29604 10265 29649
rect 10119 29558 10169 29604
rect 10215 29558 10265 29604
rect 10119 29286 10265 29558
rect 10119 29240 10169 29286
rect 10215 29240 10265 29286
rect 10119 29194 10265 29240
rect 10738 29604 10884 29649
rect 10738 29558 10788 29604
rect 10834 29558 10884 29604
rect 10738 29286 10884 29558
rect 10738 29240 10788 29286
rect 10834 29240 10884 29286
rect 10738 29194 10884 29240
rect 11357 29604 11503 29649
rect 11357 29558 11407 29604
rect 11453 29558 11503 29604
rect 11357 29286 11503 29558
rect 11357 29240 11407 29286
rect 11453 29240 11503 29286
rect 11357 29194 11503 29240
rect 11976 29604 12122 29649
rect 11976 29558 12026 29604
rect 12072 29558 12122 29604
rect 11976 29286 12122 29558
rect 11976 29240 12026 29286
rect 12072 29240 12122 29286
rect 11976 29194 12122 29240
rect 12595 29604 12741 29649
rect 12595 29558 12645 29604
rect 12691 29558 12741 29604
rect 12595 29286 12741 29558
rect 12595 29240 12645 29286
rect 12691 29240 12741 29286
rect 12595 29194 12741 29240
rect 13214 29604 13360 29649
rect 13214 29558 13264 29604
rect 13310 29558 13360 29604
rect 13214 29286 13360 29558
rect 13214 29240 13264 29286
rect 13310 29240 13360 29286
rect 13214 29194 13360 29240
rect 13833 29604 13979 29649
rect 13833 29558 13883 29604
rect 13929 29558 13979 29604
rect 13833 29286 13979 29558
rect 13833 29240 13883 29286
rect 13929 29240 13979 29286
rect 13833 29194 13979 29240
rect 14452 29604 14598 29649
rect 14452 29558 14502 29604
rect 14548 29558 14598 29604
rect 14452 29286 14598 29558
rect 14452 29240 14502 29286
rect 14548 29240 14598 29286
rect 14452 29194 14598 29240
rect 15071 29604 15217 29649
rect 15071 29558 15121 29604
rect 15167 29558 15217 29604
rect 15071 29286 15217 29558
rect 15071 29240 15121 29286
rect 15167 29240 15217 29286
rect 15071 29194 15217 29240
rect 15690 29604 15836 29649
rect 15690 29558 15740 29604
rect 15786 29558 15836 29604
rect 15690 29286 15836 29558
rect 15690 29240 15740 29286
rect 15786 29240 15836 29286
rect 15690 29194 15836 29240
rect 16309 29604 16455 29649
rect 16309 29558 16359 29604
rect 16405 29558 16455 29604
rect 16309 29286 16455 29558
rect 16309 29240 16359 29286
rect 16405 29240 16455 29286
rect 16309 29194 16455 29240
rect 16928 29604 17074 29649
rect 16928 29558 16978 29604
rect 17024 29558 17074 29604
rect 16928 29286 17074 29558
rect 16928 29240 16978 29286
rect 17024 29240 17074 29286
rect 16928 29194 17074 29240
rect 17547 29604 17693 29649
rect 17547 29558 17597 29604
rect 17643 29558 17693 29604
rect 17547 29286 17693 29558
rect 17547 29240 17597 29286
rect 17643 29240 17693 29286
rect 17547 29194 17693 29240
rect 18166 29604 18312 29649
rect 18166 29558 18216 29604
rect 18262 29558 18312 29604
rect 18166 29286 18312 29558
rect 18166 29240 18216 29286
rect 18262 29240 18312 29286
rect 18166 29194 18312 29240
rect 18785 29604 18931 29649
rect 18785 29558 18835 29604
rect 18881 29558 18931 29604
rect 18785 29286 18931 29558
rect 18785 29240 18835 29286
rect 18881 29240 18931 29286
rect 18785 29194 18931 29240
rect 19404 29604 19550 29649
rect 19404 29558 19454 29604
rect 19500 29558 19550 29604
rect 19404 29286 19550 29558
rect 19404 29240 19454 29286
rect 19500 29240 19550 29286
rect 19404 29194 19550 29240
rect 20023 29604 20169 29649
rect 20023 29558 20073 29604
rect 20119 29558 20169 29604
rect 20023 29286 20169 29558
rect 20023 29240 20073 29286
rect 20119 29240 20169 29286
rect 20023 29194 20169 29240
rect 20642 29604 20788 29649
rect 20642 29558 20692 29604
rect 20738 29558 20788 29604
rect 20642 29286 20788 29558
rect 20642 29240 20692 29286
rect 20738 29240 20788 29286
rect 20642 29194 20788 29240
rect 21261 29604 21407 29649
rect 21261 29558 21311 29604
rect 21357 29558 21407 29604
rect 21261 29286 21407 29558
rect 21261 29240 21311 29286
rect 21357 29240 21407 29286
rect 21261 29194 21407 29240
rect 21880 29604 22026 29649
rect 21880 29558 21930 29604
rect 21976 29558 22026 29604
rect 21880 29286 22026 29558
rect 21880 29240 21930 29286
rect 21976 29240 22026 29286
rect 21880 29194 22026 29240
rect 22499 29604 22639 29649
rect 22499 29558 22549 29604
rect 22595 29558 22639 29604
rect 22499 29286 22639 29558
rect 22499 29240 22549 29286
rect 22595 29240 22639 29286
rect 22499 29194 22639 29240
rect 23052 28587 23220 28632
rect 23052 28541 23143 28587
rect 23189 28541 23220 28587
rect 23052 28405 23220 28541
rect 23052 28359 23143 28405
rect 23189 28359 23220 28405
rect 23052 28224 23220 28359
rect 23052 28178 23143 28224
rect 23189 28178 23220 28224
rect 23052 28042 23220 28178
rect 23052 27996 23143 28042
rect 23189 27996 23220 28042
rect 23052 27950 23220 27996
rect 23340 28587 23444 28632
rect 23340 28541 23369 28587
rect 23415 28541 23444 28587
rect 23340 28405 23444 28541
rect 23340 28359 23369 28405
rect 23415 28359 23444 28405
rect 23340 28224 23444 28359
rect 23340 28178 23369 28224
rect 23415 28178 23444 28224
rect 23340 28042 23444 28178
rect 23340 27996 23369 28042
rect 23415 27996 23444 28042
rect 23340 27950 23444 27996
rect 23564 28587 23769 28632
rect 23564 28541 23679 28587
rect 23725 28541 23769 28587
rect 23564 28405 23769 28541
rect 23564 28359 23679 28405
rect 23725 28359 23769 28405
rect 23564 28224 23769 28359
rect 23564 28178 23679 28224
rect 23725 28178 23769 28224
rect 23564 28042 23769 28178
rect 23564 27996 23679 28042
rect 23725 27996 23769 28042
rect 23564 27950 23769 27996
rect 23052 27811 23220 27857
rect 23052 27765 23143 27811
rect 23189 27765 23220 27811
rect 23052 27630 23220 27765
rect 23052 27584 23143 27630
rect 23189 27584 23220 27630
rect 23052 27449 23220 27584
rect 23052 27403 23143 27449
rect 23189 27403 23220 27449
rect 23052 27267 23220 27403
rect 23052 27221 23143 27267
rect 23189 27221 23220 27267
rect 23052 27175 23220 27221
rect 23340 27811 23444 27857
rect 23340 27765 23369 27811
rect 23415 27765 23444 27811
rect 23340 27630 23444 27765
rect 23340 27584 23369 27630
rect 23415 27584 23444 27630
rect 23340 27449 23444 27584
rect 23340 27403 23369 27449
rect 23415 27403 23444 27449
rect 23340 27267 23444 27403
rect 23340 27221 23369 27267
rect 23415 27221 23444 27267
rect 23340 27175 23444 27221
rect 23564 27811 23769 27857
rect 23564 27765 23679 27811
rect 23725 27765 23769 27811
rect 23564 27630 23769 27765
rect 23564 27584 23679 27630
rect 23725 27584 23769 27630
rect 23564 27449 23769 27584
rect 23564 27403 23679 27449
rect 23725 27403 23769 27449
rect 23564 27267 23769 27403
rect 23564 27221 23679 27267
rect 23725 27221 23769 27267
rect 23564 27175 23769 27221
rect 23246 26943 23334 26956
rect 23246 26897 23259 26943
rect 23305 26897 23334 26943
rect 23246 26835 23334 26897
rect 23246 26789 23259 26835
rect 23305 26789 23334 26835
rect 23246 26727 23334 26789
rect 23246 26681 23259 26727
rect 23305 26681 23334 26727
rect 23246 26619 23334 26681
rect 23246 26573 23259 26619
rect 23305 26573 23334 26619
rect 23246 26511 23334 26573
rect 23246 26465 23259 26511
rect 23305 26465 23334 26511
rect 23246 26403 23334 26465
rect 23246 26357 23259 26403
rect 23305 26357 23334 26403
rect 23246 26295 23334 26357
rect 23246 26249 23259 26295
rect 23305 26249 23334 26295
rect 23246 26188 23334 26249
rect 23246 26142 23259 26188
rect 23305 26142 23334 26188
rect 23246 26081 23334 26142
rect 23246 26035 23259 26081
rect 23305 26035 23334 26081
rect 23246 25974 23334 26035
rect 23246 25928 23259 25974
rect 23305 25928 23334 25974
rect 23246 25867 23334 25928
rect 23246 25821 23259 25867
rect 23305 25821 23334 25867
rect 23246 25760 23334 25821
rect 23246 25714 23259 25760
rect 23305 25714 23334 25760
rect 23246 25653 23334 25714
rect 23246 25607 23259 25653
rect 23305 25607 23334 25653
rect 23246 25594 23334 25607
rect 23454 26943 23542 26956
rect 23454 26897 23483 26943
rect 23529 26897 23542 26943
rect 23454 26835 23542 26897
rect 23454 26789 23483 26835
rect 23529 26789 23542 26835
rect 23454 26727 23542 26789
rect 23454 26681 23483 26727
rect 23529 26681 23542 26727
rect 23454 26619 23542 26681
rect 23454 26573 23483 26619
rect 23529 26573 23542 26619
rect 23454 26511 23542 26573
rect 23454 26465 23483 26511
rect 23529 26465 23542 26511
rect 23454 26403 23542 26465
rect 23454 26357 23483 26403
rect 23529 26357 23542 26403
rect 23454 26295 23542 26357
rect 23454 26249 23483 26295
rect 23529 26249 23542 26295
rect 23454 26188 23542 26249
rect 23454 26142 23483 26188
rect 23529 26142 23542 26188
rect 23454 26081 23542 26142
rect 23454 26035 23483 26081
rect 23529 26035 23542 26081
rect 23454 25974 23542 26035
rect 23454 25928 23483 25974
rect 23529 25928 23542 25974
rect 23454 25867 23542 25928
rect 23454 25821 23483 25867
rect 23529 25821 23542 25867
rect 23454 25760 23542 25821
rect 23454 25714 23483 25760
rect 23529 25714 23542 25760
rect 23454 25653 23542 25714
rect 23454 25607 23483 25653
rect 23529 25607 23542 25653
rect 23454 25594 23542 25607
rect 23244 25356 23332 25369
rect 23244 25310 23257 25356
rect 23303 25310 23332 25356
rect 23244 25248 23332 25310
rect 23244 25202 23257 25248
rect 23303 25202 23332 25248
rect 23244 25140 23332 25202
rect 23244 25094 23257 25140
rect 23303 25094 23332 25140
rect 23244 25032 23332 25094
rect 23244 24986 23257 25032
rect 23303 24986 23332 25032
rect 23244 24924 23332 24986
rect 23244 24878 23257 24924
rect 23303 24878 23332 24924
rect 23244 24816 23332 24878
rect 23244 24770 23257 24816
rect 23303 24770 23332 24816
rect 23244 24708 23332 24770
rect 23244 24662 23257 24708
rect 23303 24662 23332 24708
rect 23244 24601 23332 24662
rect 23244 24555 23257 24601
rect 23303 24555 23332 24601
rect 23244 24494 23332 24555
rect 23244 24448 23257 24494
rect 23303 24448 23332 24494
rect 23244 24387 23332 24448
rect 23244 24341 23257 24387
rect 23303 24341 23332 24387
rect 23244 24280 23332 24341
rect 23244 24234 23257 24280
rect 23303 24234 23332 24280
rect 23244 24173 23332 24234
rect 23244 24127 23257 24173
rect 23303 24127 23332 24173
rect 23244 24066 23332 24127
rect 23244 24020 23257 24066
rect 23303 24020 23332 24066
rect 23244 24007 23332 24020
rect 23452 25356 23540 25369
rect 23452 25310 23481 25356
rect 23527 25310 23540 25356
rect 23452 25248 23540 25310
rect 23452 25202 23481 25248
rect 23527 25202 23540 25248
rect 23452 25140 23540 25202
rect 23452 25094 23481 25140
rect 23527 25094 23540 25140
rect 23452 25032 23540 25094
rect 23452 24986 23481 25032
rect 23527 24986 23540 25032
rect 23452 24924 23540 24986
rect 23452 24878 23481 24924
rect 23527 24878 23540 24924
rect 23452 24816 23540 24878
rect 23452 24770 23481 24816
rect 23527 24770 23540 24816
rect 23452 24708 23540 24770
rect 23452 24662 23481 24708
rect 23527 24662 23540 24708
rect 23452 24601 23540 24662
rect 23452 24555 23481 24601
rect 23527 24555 23540 24601
rect 23452 24494 23540 24555
rect 23452 24448 23481 24494
rect 23527 24448 23540 24494
rect 23452 24387 23540 24448
rect 23452 24341 23481 24387
rect 23527 24341 23540 24387
rect 23452 24280 23540 24341
rect 23452 24234 23481 24280
rect 23527 24234 23540 24280
rect 23452 24173 23540 24234
rect 23452 24127 23481 24173
rect 23527 24127 23540 24173
rect 23452 24066 23540 24127
rect 23452 24020 23481 24066
rect 23527 24020 23540 24066
rect 23452 24007 23540 24020
rect 23244 19806 23332 19819
rect 23244 19760 23257 19806
rect 23303 19760 23332 19806
rect 23244 19698 23332 19760
rect 23244 19652 23257 19698
rect 23303 19652 23332 19698
rect 23244 19590 23332 19652
rect 23244 19544 23257 19590
rect 23303 19544 23332 19590
rect 23244 19482 23332 19544
rect 23244 19436 23257 19482
rect 23303 19436 23332 19482
rect 23244 19374 23332 19436
rect 23244 19328 23257 19374
rect 23303 19328 23332 19374
rect 23244 19266 23332 19328
rect 23244 19220 23257 19266
rect 23303 19220 23332 19266
rect 23244 19158 23332 19220
rect 23244 19112 23257 19158
rect 23303 19112 23332 19158
rect 23244 19051 23332 19112
rect 23244 19005 23257 19051
rect 23303 19005 23332 19051
rect 23244 18944 23332 19005
rect 23244 18898 23257 18944
rect 23303 18898 23332 18944
rect 23244 18837 23332 18898
rect 23244 18791 23257 18837
rect 23303 18791 23332 18837
rect 23244 18730 23332 18791
rect 23244 18684 23257 18730
rect 23303 18684 23332 18730
rect 23244 18623 23332 18684
rect 23244 18577 23257 18623
rect 23303 18577 23332 18623
rect 23244 18516 23332 18577
rect 23244 18470 23257 18516
rect 23303 18470 23332 18516
rect 23244 18457 23332 18470
rect 23452 19806 23540 19819
rect 23452 19760 23481 19806
rect 23527 19760 23540 19806
rect 23452 19698 23540 19760
rect 23452 19652 23481 19698
rect 23527 19652 23540 19698
rect 23452 19590 23540 19652
rect 23452 19544 23481 19590
rect 23527 19544 23540 19590
rect 23452 19482 23540 19544
rect 23452 19436 23481 19482
rect 23527 19436 23540 19482
rect 23452 19374 23540 19436
rect 23452 19328 23481 19374
rect 23527 19328 23540 19374
rect 23452 19266 23540 19328
rect 23452 19220 23481 19266
rect 23527 19220 23540 19266
rect 23452 19158 23540 19220
rect 23452 19112 23481 19158
rect 23527 19112 23540 19158
rect 23452 19051 23540 19112
rect 23452 19005 23481 19051
rect 23527 19005 23540 19051
rect 23452 18944 23540 19005
rect 23452 18898 23481 18944
rect 23527 18898 23540 18944
rect 23452 18837 23540 18898
rect 23452 18791 23481 18837
rect 23527 18791 23540 18837
rect 23452 18730 23540 18791
rect 23452 18684 23481 18730
rect 23527 18684 23540 18730
rect 23452 18623 23540 18684
rect 23452 18577 23481 18623
rect 23527 18577 23540 18623
rect 23452 18516 23540 18577
rect 23452 18470 23481 18516
rect 23527 18470 23540 18516
rect 23452 18457 23540 18470
rect 23082 17719 23263 17844
rect 23082 17673 23176 17719
rect 23222 17673 23263 17719
rect 23082 17547 23263 17673
rect 23383 17719 23515 17844
rect 23383 17673 23426 17719
rect 23472 17673 23515 17719
rect 23383 17547 23515 17673
rect 23635 17719 23769 17844
rect 23635 17673 23679 17719
rect 23725 17673 23769 17719
rect 23635 17547 23769 17673
rect 23155 15158 23243 15171
rect 23155 15112 23168 15158
rect 23214 15112 23243 15158
rect 23155 15053 23243 15112
rect 23155 15007 23168 15053
rect 23214 15007 23243 15053
rect 23155 14948 23243 15007
rect 23155 14902 23168 14948
rect 23214 14902 23243 14948
rect 23155 14843 23243 14902
rect 23155 14797 23168 14843
rect 23214 14797 23243 14843
rect 23155 14738 23243 14797
rect 23155 14692 23168 14738
rect 23214 14692 23243 14738
rect 23155 14633 23243 14692
rect 23155 14587 23168 14633
rect 23214 14587 23243 14633
rect 23155 14528 23243 14587
rect 23155 14482 23168 14528
rect 23214 14482 23243 14528
rect 23155 14469 23243 14482
rect 23363 15158 23467 15171
rect 23363 15112 23392 15158
rect 23438 15112 23467 15158
rect 23363 15053 23467 15112
rect 23363 15007 23392 15053
rect 23438 15007 23467 15053
rect 23363 14948 23467 15007
rect 23363 14902 23392 14948
rect 23438 14902 23467 14948
rect 23363 14843 23467 14902
rect 23363 14797 23392 14843
rect 23438 14797 23467 14843
rect 23363 14738 23467 14797
rect 23363 14692 23392 14738
rect 23438 14692 23467 14738
rect 23363 14633 23467 14692
rect 23363 14587 23392 14633
rect 23438 14587 23467 14633
rect 23363 14528 23467 14587
rect 23363 14482 23392 14528
rect 23438 14482 23467 14528
rect 23363 14469 23467 14482
rect 23587 15158 23675 15171
rect 23587 15112 23616 15158
rect 23662 15112 23675 15158
rect 23587 15053 23675 15112
rect 23587 15007 23616 15053
rect 23662 15007 23675 15053
rect 23587 14948 23675 15007
rect 23587 14902 23616 14948
rect 23662 14902 23675 14948
rect 23587 14843 23675 14902
rect 23587 14797 23616 14843
rect 23662 14797 23675 14843
rect 23587 14738 23675 14797
rect 23587 14692 23616 14738
rect 23662 14692 23675 14738
rect 23587 14633 23675 14692
rect 23587 14587 23616 14633
rect 23662 14587 23675 14633
rect 23587 14528 23675 14587
rect 23587 14482 23616 14528
rect 23662 14482 23675 14528
rect 23587 14469 23675 14482
rect 23159 10510 23247 10523
rect 23159 10464 23172 10510
rect 23218 10464 23247 10510
rect 23159 10407 23247 10464
rect 23159 10361 23172 10407
rect 23218 10361 23247 10407
rect 23159 10304 23247 10361
rect 23159 10258 23172 10304
rect 23218 10258 23247 10304
rect 23159 10201 23247 10258
rect 23159 10155 23172 10201
rect 23218 10155 23247 10201
rect 23159 10098 23247 10155
rect 23159 10052 23172 10098
rect 23218 10052 23247 10098
rect 23159 9995 23247 10052
rect 23159 9949 23172 9995
rect 23218 9949 23247 9995
rect 23159 9892 23247 9949
rect 23159 9846 23172 9892
rect 23218 9846 23247 9892
rect 23159 9789 23247 9846
rect 23159 9743 23172 9789
rect 23218 9743 23247 9789
rect 23159 9686 23247 9743
rect 23159 9640 23172 9686
rect 23218 9640 23247 9686
rect 23159 9583 23247 9640
rect 23159 9537 23172 9583
rect 23218 9537 23247 9583
rect 23159 9480 23247 9537
rect 23159 9434 23172 9480
rect 23218 9434 23247 9480
rect 23159 9377 23247 9434
rect 23159 9331 23172 9377
rect 23218 9331 23247 9377
rect 23159 9274 23247 9331
rect 23159 9228 23172 9274
rect 23218 9228 23247 9274
rect 23159 9171 23247 9228
rect 23159 9125 23172 9171
rect 23218 9125 23247 9171
rect 23159 9068 23247 9125
rect 23159 9022 23172 9068
rect 23218 9022 23247 9068
rect 23159 8965 23247 9022
rect 23159 8919 23172 8965
rect 23218 8919 23247 8965
rect 23159 8862 23247 8919
rect 23159 8408 23172 8862
rect 23218 8408 23247 8862
rect 23159 8395 23247 8408
rect 23367 10510 23471 10523
rect 23367 10464 23396 10510
rect 23442 10464 23471 10510
rect 23367 10407 23471 10464
rect 23367 10361 23396 10407
rect 23442 10361 23471 10407
rect 23367 10304 23471 10361
rect 23367 10258 23396 10304
rect 23442 10258 23471 10304
rect 23367 10201 23471 10258
rect 23367 10155 23396 10201
rect 23442 10155 23471 10201
rect 23367 10098 23471 10155
rect 23367 10052 23396 10098
rect 23442 10052 23471 10098
rect 23367 9995 23471 10052
rect 23367 9949 23396 9995
rect 23442 9949 23471 9995
rect 23367 9892 23471 9949
rect 23367 9846 23396 9892
rect 23442 9846 23471 9892
rect 23367 9789 23471 9846
rect 23367 9743 23396 9789
rect 23442 9743 23471 9789
rect 23367 9686 23471 9743
rect 23367 9640 23396 9686
rect 23442 9640 23471 9686
rect 23367 9583 23471 9640
rect 23367 9537 23396 9583
rect 23442 9537 23471 9583
rect 23367 9480 23471 9537
rect 23367 9434 23396 9480
rect 23442 9434 23471 9480
rect 23367 9377 23471 9434
rect 23367 9331 23396 9377
rect 23442 9331 23471 9377
rect 23367 9274 23471 9331
rect 23367 9228 23396 9274
rect 23442 9228 23471 9274
rect 23367 9171 23471 9228
rect 23367 9125 23396 9171
rect 23442 9125 23471 9171
rect 23367 9068 23471 9125
rect 23367 9022 23396 9068
rect 23442 9022 23471 9068
rect 23367 8965 23471 9022
rect 23367 8919 23396 8965
rect 23442 8919 23471 8965
rect 23367 8862 23471 8919
rect 23367 8408 23396 8862
rect 23442 8408 23471 8862
rect 23367 8395 23471 8408
rect 23591 10510 23679 10523
rect 23591 10464 23620 10510
rect 23666 10464 23679 10510
rect 23591 10407 23679 10464
rect 23591 10361 23620 10407
rect 23666 10361 23679 10407
rect 23591 10304 23679 10361
rect 23591 10258 23620 10304
rect 23666 10258 23679 10304
rect 23591 10201 23679 10258
rect 23591 10155 23620 10201
rect 23666 10155 23679 10201
rect 23591 10098 23679 10155
rect 23591 10052 23620 10098
rect 23666 10052 23679 10098
rect 23591 9995 23679 10052
rect 23591 9949 23620 9995
rect 23666 9949 23679 9995
rect 23591 9892 23679 9949
rect 23591 9846 23620 9892
rect 23666 9846 23679 9892
rect 23591 9789 23679 9846
rect 23591 9743 23620 9789
rect 23666 9743 23679 9789
rect 23591 9686 23679 9743
rect 23591 9640 23620 9686
rect 23666 9640 23679 9686
rect 23591 9583 23679 9640
rect 23591 9537 23620 9583
rect 23666 9537 23679 9583
rect 23591 9480 23679 9537
rect 23591 9434 23620 9480
rect 23666 9434 23679 9480
rect 23591 9377 23679 9434
rect 23591 9331 23620 9377
rect 23666 9331 23679 9377
rect 23591 9274 23679 9331
rect 23591 9228 23620 9274
rect 23666 9228 23679 9274
rect 23591 9171 23679 9228
rect 23591 9125 23620 9171
rect 23666 9125 23679 9171
rect 23591 9068 23679 9125
rect 23591 9022 23620 9068
rect 23666 9022 23679 9068
rect 23591 8965 23679 9022
rect 23591 8919 23620 8965
rect 23666 8919 23679 8965
rect 23591 8862 23679 8919
rect 23591 8408 23620 8862
rect 23666 8408 23679 8862
rect 23591 8395 23679 8408
<< mvndiffc >>
rect 23257 23619 23303 23665
rect 23257 23511 23303 23557
rect 23257 23403 23303 23449
rect 23257 23295 23303 23341
rect 23257 23187 23303 23233
rect 23257 23079 23303 23125
rect 23257 22971 23303 23017
rect 23257 22864 23303 22910
rect 23257 22757 23303 22803
rect 23257 22650 23303 22696
rect 23257 22543 23303 22589
rect 23257 22436 23303 22482
rect 23257 22329 23303 22375
rect 23481 23619 23527 23665
rect 23481 23511 23527 23557
rect 23481 23403 23527 23449
rect 23481 23295 23527 23341
rect 23481 23187 23527 23233
rect 23481 23079 23527 23125
rect 23481 22971 23527 23017
rect 23481 22864 23527 22910
rect 23481 22757 23527 22803
rect 23481 22650 23527 22696
rect 23481 22543 23527 22589
rect 23481 22436 23527 22482
rect 23481 22329 23527 22375
rect 23257 21615 23303 21661
rect 23257 21507 23303 21553
rect 23257 21399 23303 21445
rect 23257 21291 23303 21337
rect 23257 21183 23303 21229
rect 23257 21075 23303 21121
rect 23257 20967 23303 21013
rect 23257 20860 23303 20906
rect 23257 20753 23303 20799
rect 23257 20646 23303 20692
rect 23257 20539 23303 20585
rect 23257 20432 23303 20478
rect 23257 20325 23303 20371
rect 23481 21615 23527 21661
rect 23481 21507 23527 21553
rect 23481 21399 23527 21445
rect 23481 21291 23527 21337
rect 23481 21183 23527 21229
rect 23481 21075 23527 21121
rect 23481 20967 23527 21013
rect 23481 20860 23527 20906
rect 23481 20753 23527 20799
rect 23481 20646 23527 20692
rect 23481 20539 23527 20585
rect 23481 20432 23527 20478
rect 23481 20325 23527 20371
rect 23217 17176 23263 17222
rect 23441 17176 23487 17222
rect 23665 17176 23711 17222
rect 23168 13902 23214 14152
rect 23392 13902 23438 14152
rect 23616 13902 23662 14152
rect 23172 10817 23218 12491
rect 23396 10817 23442 12491
rect 23620 10817 23666 12491
<< mvpdiffc >>
rect 265 29558 311 29604
rect 265 29240 311 29286
rect 884 29558 930 29604
rect 884 29240 930 29286
rect 1503 29558 1549 29604
rect 1503 29240 1549 29286
rect 2122 29558 2168 29604
rect 2122 29240 2168 29286
rect 2741 29558 2787 29604
rect 2741 29240 2787 29286
rect 3360 29558 3406 29604
rect 3360 29240 3406 29286
rect 3979 29558 4025 29604
rect 3979 29240 4025 29286
rect 4598 29558 4644 29604
rect 4598 29240 4644 29286
rect 5217 29558 5263 29604
rect 5217 29240 5263 29286
rect 5836 29558 5882 29604
rect 5836 29240 5882 29286
rect 6455 29558 6501 29604
rect 6455 29240 6501 29286
rect 7074 29558 7120 29604
rect 7074 29240 7120 29286
rect 7693 29558 7739 29604
rect 7693 29240 7739 29286
rect 8312 29558 8358 29604
rect 8312 29240 8358 29286
rect 8931 29558 8977 29604
rect 8931 29240 8977 29286
rect 9550 29558 9596 29604
rect 9550 29240 9596 29286
rect 10169 29558 10215 29604
rect 10169 29240 10215 29286
rect 10788 29558 10834 29604
rect 10788 29240 10834 29286
rect 11407 29558 11453 29604
rect 11407 29240 11453 29286
rect 12026 29558 12072 29604
rect 12026 29240 12072 29286
rect 12645 29558 12691 29604
rect 12645 29240 12691 29286
rect 13264 29558 13310 29604
rect 13264 29240 13310 29286
rect 13883 29558 13929 29604
rect 13883 29240 13929 29286
rect 14502 29558 14548 29604
rect 14502 29240 14548 29286
rect 15121 29558 15167 29604
rect 15121 29240 15167 29286
rect 15740 29558 15786 29604
rect 15740 29240 15786 29286
rect 16359 29558 16405 29604
rect 16359 29240 16405 29286
rect 16978 29558 17024 29604
rect 16978 29240 17024 29286
rect 17597 29558 17643 29604
rect 17597 29240 17643 29286
rect 18216 29558 18262 29604
rect 18216 29240 18262 29286
rect 18835 29558 18881 29604
rect 18835 29240 18881 29286
rect 19454 29558 19500 29604
rect 19454 29240 19500 29286
rect 20073 29558 20119 29604
rect 20073 29240 20119 29286
rect 20692 29558 20738 29604
rect 20692 29240 20738 29286
rect 21311 29558 21357 29604
rect 21311 29240 21357 29286
rect 21930 29558 21976 29604
rect 21930 29240 21976 29286
rect 22549 29558 22595 29604
rect 22549 29240 22595 29286
rect 23143 28541 23189 28587
rect 23143 28359 23189 28405
rect 23143 28178 23189 28224
rect 23143 27996 23189 28042
rect 23369 28541 23415 28587
rect 23369 28359 23415 28405
rect 23369 28178 23415 28224
rect 23369 27996 23415 28042
rect 23679 28541 23725 28587
rect 23679 28359 23725 28405
rect 23679 28178 23725 28224
rect 23679 27996 23725 28042
rect 23143 27765 23189 27811
rect 23143 27584 23189 27630
rect 23143 27403 23189 27449
rect 23143 27221 23189 27267
rect 23369 27765 23415 27811
rect 23369 27584 23415 27630
rect 23369 27403 23415 27449
rect 23369 27221 23415 27267
rect 23679 27765 23725 27811
rect 23679 27584 23725 27630
rect 23679 27403 23725 27449
rect 23679 27221 23725 27267
rect 23259 26897 23305 26943
rect 23259 26789 23305 26835
rect 23259 26681 23305 26727
rect 23259 26573 23305 26619
rect 23259 26465 23305 26511
rect 23259 26357 23305 26403
rect 23259 26249 23305 26295
rect 23259 26142 23305 26188
rect 23259 26035 23305 26081
rect 23259 25928 23305 25974
rect 23259 25821 23305 25867
rect 23259 25714 23305 25760
rect 23259 25607 23305 25653
rect 23483 26897 23529 26943
rect 23483 26789 23529 26835
rect 23483 26681 23529 26727
rect 23483 26573 23529 26619
rect 23483 26465 23529 26511
rect 23483 26357 23529 26403
rect 23483 26249 23529 26295
rect 23483 26142 23529 26188
rect 23483 26035 23529 26081
rect 23483 25928 23529 25974
rect 23483 25821 23529 25867
rect 23483 25714 23529 25760
rect 23483 25607 23529 25653
rect 23257 25310 23303 25356
rect 23257 25202 23303 25248
rect 23257 25094 23303 25140
rect 23257 24986 23303 25032
rect 23257 24878 23303 24924
rect 23257 24770 23303 24816
rect 23257 24662 23303 24708
rect 23257 24555 23303 24601
rect 23257 24448 23303 24494
rect 23257 24341 23303 24387
rect 23257 24234 23303 24280
rect 23257 24127 23303 24173
rect 23257 24020 23303 24066
rect 23481 25310 23527 25356
rect 23481 25202 23527 25248
rect 23481 25094 23527 25140
rect 23481 24986 23527 25032
rect 23481 24878 23527 24924
rect 23481 24770 23527 24816
rect 23481 24662 23527 24708
rect 23481 24555 23527 24601
rect 23481 24448 23527 24494
rect 23481 24341 23527 24387
rect 23481 24234 23527 24280
rect 23481 24127 23527 24173
rect 23481 24020 23527 24066
rect 23257 19760 23303 19806
rect 23257 19652 23303 19698
rect 23257 19544 23303 19590
rect 23257 19436 23303 19482
rect 23257 19328 23303 19374
rect 23257 19220 23303 19266
rect 23257 19112 23303 19158
rect 23257 19005 23303 19051
rect 23257 18898 23303 18944
rect 23257 18791 23303 18837
rect 23257 18684 23303 18730
rect 23257 18577 23303 18623
rect 23257 18470 23303 18516
rect 23481 19760 23527 19806
rect 23481 19652 23527 19698
rect 23481 19544 23527 19590
rect 23481 19436 23527 19482
rect 23481 19328 23527 19374
rect 23481 19220 23527 19266
rect 23481 19112 23527 19158
rect 23481 19005 23527 19051
rect 23481 18898 23527 18944
rect 23481 18791 23527 18837
rect 23481 18684 23527 18730
rect 23481 18577 23527 18623
rect 23481 18470 23527 18516
rect 23176 17673 23222 17719
rect 23426 17673 23472 17719
rect 23679 17673 23725 17719
rect 23168 15112 23214 15158
rect 23168 15007 23214 15053
rect 23168 14902 23214 14948
rect 23168 14797 23214 14843
rect 23168 14692 23214 14738
rect 23168 14587 23214 14633
rect 23168 14482 23214 14528
rect 23392 15112 23438 15158
rect 23392 15007 23438 15053
rect 23392 14902 23438 14948
rect 23392 14797 23438 14843
rect 23392 14692 23438 14738
rect 23392 14587 23438 14633
rect 23392 14482 23438 14528
rect 23616 15112 23662 15158
rect 23616 15007 23662 15053
rect 23616 14902 23662 14948
rect 23616 14797 23662 14843
rect 23616 14692 23662 14738
rect 23616 14587 23662 14633
rect 23616 14482 23662 14528
rect 23172 10464 23218 10510
rect 23172 10361 23218 10407
rect 23172 10258 23218 10304
rect 23172 10155 23218 10201
rect 23172 10052 23218 10098
rect 23172 9949 23218 9995
rect 23172 9846 23218 9892
rect 23172 9743 23218 9789
rect 23172 9640 23218 9686
rect 23172 9537 23218 9583
rect 23172 9434 23218 9480
rect 23172 9331 23218 9377
rect 23172 9228 23218 9274
rect 23172 9125 23218 9171
rect 23172 9022 23218 9068
rect 23172 8919 23218 8965
rect 23172 8408 23218 8862
rect 23396 10464 23442 10510
rect 23396 10361 23442 10407
rect 23396 10258 23442 10304
rect 23396 10155 23442 10201
rect 23396 10052 23442 10098
rect 23396 9949 23442 9995
rect 23396 9846 23442 9892
rect 23396 9743 23442 9789
rect 23396 9640 23442 9686
rect 23396 9537 23442 9583
rect 23396 9434 23442 9480
rect 23396 9331 23442 9377
rect 23396 9228 23442 9274
rect 23396 9125 23442 9171
rect 23396 9022 23442 9068
rect 23396 8919 23442 8965
rect 23396 8408 23442 8862
rect 23620 10464 23666 10510
rect 23620 10361 23666 10407
rect 23620 10258 23666 10304
rect 23620 10155 23666 10201
rect 23620 10052 23666 10098
rect 23620 9949 23666 9995
rect 23620 9846 23666 9892
rect 23620 9743 23666 9789
rect 23620 9640 23666 9686
rect 23620 9537 23666 9583
rect 23620 9434 23666 9480
rect 23620 9331 23666 9377
rect 23620 9228 23666 9274
rect 23620 9125 23666 9171
rect 23620 9022 23666 9068
rect 23620 8919 23666 8965
rect 23620 8408 23666 8862
<< mvpsubdiff >>
rect 23622 22019 23782 22079
rect 23622 21973 23679 22019
rect 23725 21973 23782 22019
rect 23622 21913 23782 21973
rect 23228 16923 23688 16942
rect 23228 16877 23247 16923
rect 23669 16877 23688 16923
rect 23228 16858 23688 16877
rect 23176 13613 23652 13673
rect 23176 13567 23233 13613
rect 23279 13567 23391 13613
rect 23437 13567 23549 13613
rect 23595 13567 23652 13613
rect 23176 13507 23652 13567
<< mvnsubdiff >>
rect 23052 28924 23703 28981
rect 23052 28878 23211 28924
rect 23257 28878 23369 28924
rect 23415 28878 23527 28924
rect 23573 28878 23703 28924
rect 23052 28821 23703 28878
rect 23082 18174 23780 18231
rect 23082 18128 23205 18174
rect 23251 18128 23363 18174
rect 23409 18128 23521 18174
rect 23567 18128 23679 18174
rect 23725 18128 23780 18174
rect 23082 18071 23780 18128
rect 23121 15608 23593 15665
rect 23121 15562 23176 15608
rect 23222 15562 23334 15608
rect 23380 15562 23492 15608
rect 23538 15562 23593 15608
rect 23121 15505 23593 15562
rect 23004 7288 23159 7345
rect 23004 7242 23058 7288
rect 23104 7242 23159 7288
rect 23004 7185 23159 7242
rect 23548 7288 23703 7345
rect 23548 7242 23602 7288
rect 23648 7242 23703 7288
rect 23548 7185 23703 7242
<< mvpsubdiffcont >>
rect 23679 21973 23725 22019
rect 23247 16877 23669 16923
rect 23233 13567 23279 13613
rect 23391 13567 23437 13613
rect 23549 13567 23595 13613
<< mvnsubdiffcont >>
rect 23211 28878 23257 28924
rect 23369 28878 23415 28924
rect 23527 28878 23573 28924
rect 23205 18128 23251 18174
rect 23363 18128 23409 18174
rect 23521 18128 23567 18174
rect 23679 18128 23725 18174
rect 23176 15562 23222 15608
rect 23334 15562 23380 15608
rect 23492 15562 23538 15608
rect 23058 7242 23104 7288
rect 23602 7242 23648 7288
<< polysilicon >>
rect 50 89536 364 89555
rect 50 89396 69 89536
rect 115 89401 364 89536
rect 23648 89472 24018 89555
rect 23648 89426 23899 89472
rect 23945 89426 24018 89472
rect 23648 89401 24018 89426
rect 115 89396 134 89401
rect 50 89377 134 89396
rect 23826 89308 24018 89401
rect 23826 89262 23899 89308
rect 23945 89262 24018 89308
rect 23826 89216 24018 89262
rect 50 87877 364 88013
rect 50 87737 69 87877
rect 115 87859 364 87877
rect 23648 87912 24018 88013
rect 23648 87866 23899 87912
rect 23945 87866 24018 87912
rect 23648 87859 24018 87866
rect 115 87755 134 87859
rect 23826 87755 24018 87859
rect 115 87737 364 87755
rect 50 87601 364 87737
rect 23648 87748 24018 87755
rect 23648 87702 23899 87748
rect 23945 87702 24018 87748
rect 23648 87601 24018 87702
rect 50 86077 364 86213
rect 50 85937 69 86077
rect 115 86059 364 86077
rect 23648 86112 24018 86213
rect 23648 86066 23899 86112
rect 23945 86066 24018 86112
rect 23648 86059 24018 86066
rect 115 85955 134 86059
rect 23826 85955 24018 86059
rect 115 85937 364 85955
rect 50 85801 364 85937
rect 23648 85948 24018 85955
rect 23648 85902 23899 85948
rect 23945 85902 24018 85948
rect 23648 85801 24018 85902
rect 50 84277 364 84413
rect 50 84137 69 84277
rect 115 84259 364 84277
rect 23648 84312 24018 84413
rect 23648 84266 23899 84312
rect 23945 84266 24018 84312
rect 23648 84259 24018 84266
rect 115 84155 134 84259
rect 23826 84155 24018 84259
rect 115 84137 364 84155
rect 50 84001 364 84137
rect 23648 84148 24018 84155
rect 23648 84102 23899 84148
rect 23945 84102 24018 84148
rect 23648 84001 24018 84102
rect 50 82477 364 82613
rect 50 82337 69 82477
rect 115 82459 364 82477
rect 23648 82512 24018 82613
rect 23648 82466 23899 82512
rect 23945 82466 24018 82512
rect 23648 82459 24018 82466
rect 115 82355 134 82459
rect 23826 82355 24018 82459
rect 115 82337 364 82355
rect 50 82201 364 82337
rect 23648 82348 24018 82355
rect 23648 82302 23899 82348
rect 23945 82302 24018 82348
rect 23648 82201 24018 82302
rect 50 80677 364 80813
rect 50 80537 69 80677
rect 115 80659 364 80677
rect 23648 80712 24018 80813
rect 23648 80666 23899 80712
rect 23945 80666 24018 80712
rect 23648 80659 24018 80666
rect 115 80555 134 80659
rect 23826 80555 24018 80659
rect 115 80537 364 80555
rect 50 80401 364 80537
rect 23648 80548 24018 80555
rect 23648 80502 23899 80548
rect 23945 80502 24018 80548
rect 23648 80401 24018 80502
rect 50 78877 364 79013
rect 50 78737 69 78877
rect 115 78859 364 78877
rect 23648 78912 24018 79013
rect 23648 78866 23899 78912
rect 23945 78866 24018 78912
rect 23648 78859 24018 78866
rect 115 78755 134 78859
rect 23826 78755 24018 78859
rect 115 78737 364 78755
rect 50 78601 364 78737
rect 23648 78748 24018 78755
rect 23648 78702 23899 78748
rect 23945 78702 24018 78748
rect 23648 78601 24018 78702
rect 50 77077 364 77213
rect 50 76937 69 77077
rect 115 77059 364 77077
rect 23648 77112 24018 77213
rect 23648 77066 23899 77112
rect 23945 77066 24018 77112
rect 23648 77059 24018 77066
rect 115 76955 134 77059
rect 23826 76955 24018 77059
rect 115 76937 364 76955
rect 50 76801 364 76937
rect 23648 76948 24018 76955
rect 23648 76902 23899 76948
rect 23945 76902 24018 76948
rect 23648 76801 24018 76902
rect 50 75277 364 75413
rect 50 75137 69 75277
rect 115 75259 364 75277
rect 23648 75312 24018 75413
rect 23648 75266 23899 75312
rect 23945 75266 24018 75312
rect 23648 75259 24018 75266
rect 115 75155 134 75259
rect 23826 75155 24018 75259
rect 115 75137 364 75155
rect 50 75001 364 75137
rect 23648 75148 24018 75155
rect 23648 75102 23899 75148
rect 23945 75102 24018 75148
rect 23648 75001 24018 75102
rect 50 73477 364 73613
rect 50 73337 69 73477
rect 115 73459 364 73477
rect 23648 73512 24018 73613
rect 23648 73466 23899 73512
rect 23945 73466 24018 73512
rect 23648 73459 24018 73466
rect 115 73355 134 73459
rect 23826 73355 24018 73459
rect 115 73337 364 73355
rect 50 73201 364 73337
rect 23648 73348 24018 73355
rect 23648 73302 23899 73348
rect 23945 73302 24018 73348
rect 23648 73201 24018 73302
rect 50 71677 364 71813
rect 50 71537 69 71677
rect 115 71659 364 71677
rect 23648 71712 24018 71813
rect 23648 71666 23899 71712
rect 23945 71666 24018 71712
rect 23648 71659 24018 71666
rect 115 71555 134 71659
rect 23826 71555 24018 71659
rect 115 71537 364 71555
rect 50 71401 364 71537
rect 23648 71548 24018 71555
rect 23648 71502 23899 71548
rect 23945 71502 24018 71548
rect 23648 71401 24018 71502
rect 50 69877 364 70013
rect 50 69737 69 69877
rect 115 69859 364 69877
rect 23648 69912 24018 70013
rect 23648 69866 23899 69912
rect 23945 69866 24018 69912
rect 23648 69859 24018 69866
rect 115 69755 134 69859
rect 23826 69755 24018 69859
rect 115 69737 364 69755
rect 50 69601 364 69737
rect 23648 69748 24018 69755
rect 23648 69702 23899 69748
rect 23945 69702 24018 69748
rect 23648 69601 24018 69702
rect 50 68077 364 68213
rect 50 67937 69 68077
rect 115 68059 364 68077
rect 23648 68112 24018 68213
rect 23648 68066 23899 68112
rect 23945 68066 24018 68112
rect 23648 68059 24018 68066
rect 115 67955 134 68059
rect 23826 67955 24018 68059
rect 115 67937 364 67955
rect 50 67801 364 67937
rect 23648 67948 24018 67955
rect 23648 67902 23899 67948
rect 23945 67902 24018 67948
rect 23648 67801 24018 67902
rect 50 66277 364 66413
rect 50 66137 69 66277
rect 115 66259 364 66277
rect 23648 66312 24018 66413
rect 23648 66266 23899 66312
rect 23945 66266 24018 66312
rect 23648 66259 24018 66266
rect 115 66155 134 66259
rect 23826 66155 24018 66259
rect 115 66137 364 66155
rect 50 66001 364 66137
rect 23648 66148 24018 66155
rect 23648 66102 23899 66148
rect 23945 66102 24018 66148
rect 23648 66001 24018 66102
rect 50 64477 364 64613
rect 50 64337 69 64477
rect 115 64459 364 64477
rect 23648 64512 24018 64613
rect 23648 64466 23899 64512
rect 23945 64466 24018 64512
rect 23648 64459 24018 64466
rect 115 64355 134 64459
rect 23826 64355 24018 64459
rect 115 64337 364 64355
rect 50 64201 364 64337
rect 23648 64348 24018 64355
rect 23648 64302 23899 64348
rect 23945 64302 24018 64348
rect 23648 64201 24018 64302
rect 50 62677 364 62813
rect 50 62537 69 62677
rect 115 62659 364 62677
rect 23648 62712 24018 62813
rect 23648 62666 23899 62712
rect 23945 62666 24018 62712
rect 23648 62659 24018 62666
rect 115 62555 134 62659
rect 23826 62555 24018 62659
rect 115 62537 364 62555
rect 50 62401 364 62537
rect 23648 62548 24018 62555
rect 23648 62502 23899 62548
rect 23945 62502 24018 62548
rect 23648 62401 24018 62502
rect 50 60877 364 61013
rect 50 60737 69 60877
rect 115 60859 364 60877
rect 23648 60912 24018 61013
rect 23648 60866 23899 60912
rect 23945 60866 24018 60912
rect 23648 60859 24018 60866
rect 115 60755 134 60859
rect 23826 60755 24018 60859
rect 115 60737 364 60755
rect 50 60601 364 60737
rect 23648 60748 24018 60755
rect 23648 60702 23899 60748
rect 23945 60702 24018 60748
rect 23648 60601 24018 60702
rect 50 59077 364 59213
rect 50 58937 69 59077
rect 115 59059 364 59077
rect 23648 59112 24018 59213
rect 23648 59066 23899 59112
rect 23945 59066 24018 59112
rect 23648 59059 24018 59066
rect 115 58955 134 59059
rect 23826 58955 24018 59059
rect 115 58937 364 58955
rect 50 58801 364 58937
rect 23648 58948 24018 58955
rect 23648 58902 23899 58948
rect 23945 58902 24018 58948
rect 23648 58801 24018 58902
rect 50 57277 364 57413
rect 50 57137 69 57277
rect 115 57259 364 57277
rect 23648 57312 24018 57413
rect 23648 57266 23899 57312
rect 23945 57266 24018 57312
rect 23648 57259 24018 57266
rect 115 57155 134 57259
rect 23826 57155 24018 57259
rect 115 57137 364 57155
rect 50 57001 364 57137
rect 23648 57148 24018 57155
rect 23648 57102 23899 57148
rect 23945 57102 24018 57148
rect 23648 57001 24018 57102
rect 50 55477 364 55613
rect 50 55337 69 55477
rect 115 55459 364 55477
rect 23648 55512 24018 55613
rect 23648 55466 23899 55512
rect 23945 55466 24018 55512
rect 23648 55459 24018 55466
rect 115 55355 134 55459
rect 23826 55355 24018 55459
rect 115 55337 364 55355
rect 50 55201 364 55337
rect 23648 55348 24018 55355
rect 23648 55302 23899 55348
rect 23945 55302 24018 55348
rect 23648 55201 24018 55302
rect 50 53677 364 53813
rect 50 53537 69 53677
rect 115 53659 364 53677
rect 23648 53712 24018 53813
rect 23648 53666 23899 53712
rect 23945 53666 24018 53712
rect 23648 53659 24018 53666
rect 115 53555 134 53659
rect 23826 53555 24018 53659
rect 115 53537 364 53555
rect 50 53401 364 53537
rect 23648 53548 24018 53555
rect 23648 53502 23899 53548
rect 23945 53502 24018 53548
rect 23648 53401 24018 53502
rect 50 51877 364 52013
rect 50 51737 69 51877
rect 115 51859 364 51877
rect 23648 51912 24018 52013
rect 23648 51866 23899 51912
rect 23945 51866 24018 51912
rect 23648 51859 24018 51866
rect 115 51755 134 51859
rect 23826 51755 24018 51859
rect 115 51737 364 51755
rect 50 51601 364 51737
rect 23648 51748 24018 51755
rect 23648 51702 23899 51748
rect 23945 51702 24018 51748
rect 23648 51601 24018 51702
rect 50 50077 364 50213
rect 50 49937 69 50077
rect 115 50059 364 50077
rect 23648 50112 24018 50213
rect 23648 50066 23899 50112
rect 23945 50066 24018 50112
rect 23648 50059 24018 50066
rect 115 49955 134 50059
rect 23826 49955 24018 50059
rect 115 49937 364 49955
rect 50 49801 364 49937
rect 23648 49948 24018 49955
rect 23648 49902 23899 49948
rect 23945 49902 24018 49948
rect 23648 49801 24018 49902
rect 50 48277 364 48413
rect 50 48137 69 48277
rect 115 48259 364 48277
rect 23648 48312 24018 48413
rect 23648 48266 23899 48312
rect 23945 48266 24018 48312
rect 23648 48259 24018 48266
rect 115 48155 134 48259
rect 23826 48155 24018 48259
rect 115 48137 364 48155
rect 50 48001 364 48137
rect 23648 48148 24018 48155
rect 23648 48102 23899 48148
rect 23945 48102 24018 48148
rect 23648 48001 24018 48102
rect 50 46477 364 46613
rect 50 46337 69 46477
rect 115 46459 364 46477
rect 23648 46512 24018 46613
rect 23648 46466 23899 46512
rect 23945 46466 24018 46512
rect 23648 46459 24018 46466
rect 115 46355 134 46459
rect 23826 46355 24018 46459
rect 115 46337 364 46355
rect 50 46201 364 46337
rect 23648 46348 24018 46355
rect 23648 46302 23899 46348
rect 23945 46302 24018 46348
rect 23648 46201 24018 46302
rect 50 44677 364 44813
rect 50 44537 69 44677
rect 115 44659 364 44677
rect 23648 44712 24018 44813
rect 23648 44666 23899 44712
rect 23945 44666 24018 44712
rect 23648 44659 24018 44666
rect 115 44555 134 44659
rect 23826 44555 24018 44659
rect 115 44537 364 44555
rect 50 44401 364 44537
rect 23648 44548 24018 44555
rect 23648 44502 23899 44548
rect 23945 44502 24018 44548
rect 23648 44401 24018 44502
rect 50 42877 364 43013
rect 50 42737 69 42877
rect 115 42859 364 42877
rect 23648 42912 24018 43013
rect 23648 42866 23899 42912
rect 23945 42866 24018 42912
rect 23648 42859 24018 42866
rect 115 42755 134 42859
rect 23826 42755 24018 42859
rect 115 42737 364 42755
rect 50 42601 364 42737
rect 23648 42748 24018 42755
rect 23648 42702 23899 42748
rect 23945 42702 24018 42748
rect 23648 42601 24018 42702
rect 50 41077 364 41213
rect 50 40937 69 41077
rect 115 41059 364 41077
rect 23648 41112 24018 41213
rect 23648 41066 23899 41112
rect 23945 41066 24018 41112
rect 23648 41059 24018 41066
rect 115 40955 134 41059
rect 23826 40955 24018 41059
rect 115 40937 364 40955
rect 50 40801 364 40937
rect 23648 40948 24018 40955
rect 23648 40902 23899 40948
rect 23945 40902 24018 40948
rect 23648 40801 24018 40902
rect 50 39277 364 39413
rect 50 39137 69 39277
rect 115 39259 364 39277
rect 23648 39312 24018 39413
rect 23648 39266 23899 39312
rect 23945 39266 24018 39312
rect 23648 39259 24018 39266
rect 115 39155 134 39259
rect 23826 39155 24018 39259
rect 115 39137 364 39155
rect 50 39001 364 39137
rect 23648 39148 24018 39155
rect 23648 39102 23899 39148
rect 23945 39102 24018 39148
rect 23648 39001 24018 39102
rect 50 37477 364 37613
rect 50 37337 69 37477
rect 115 37459 364 37477
rect 23648 37512 24018 37613
rect 23648 37466 23899 37512
rect 23945 37466 24018 37512
rect 23648 37459 24018 37466
rect 115 37355 134 37459
rect 23826 37355 24018 37459
rect 115 37337 364 37355
rect 50 37201 364 37337
rect 23648 37348 24018 37355
rect 23648 37302 23899 37348
rect 23945 37302 24018 37348
rect 23648 37201 24018 37302
rect 50 35677 364 35813
rect 50 35537 69 35677
rect 115 35659 364 35677
rect 23648 35712 24018 35813
rect 23648 35666 23899 35712
rect 23945 35666 24018 35712
rect 23648 35659 24018 35666
rect 115 35555 134 35659
rect 23826 35555 24018 35659
rect 115 35537 364 35555
rect 50 35401 364 35537
rect 23648 35548 24018 35555
rect 23648 35502 23899 35548
rect 23945 35502 24018 35548
rect 23648 35401 24018 35502
rect 50 33877 364 34013
rect 50 33737 69 33877
rect 115 33859 364 33877
rect 23648 33912 24018 34013
rect 23648 33866 23899 33912
rect 23945 33866 24018 33912
rect 23648 33859 24018 33866
rect 115 33755 134 33859
rect 23826 33755 24018 33859
rect 115 33737 364 33755
rect 50 33601 364 33737
rect 23648 33748 24018 33755
rect 23648 33702 23899 33748
rect 23945 33702 24018 33748
rect 23648 33601 24018 33702
rect 50 32077 364 32213
rect 50 31937 69 32077
rect 115 32059 364 32077
rect 23648 32112 24018 32213
rect 23648 32066 23899 32112
rect 23945 32066 24018 32112
rect 23648 32059 24018 32066
rect 115 31955 134 32059
rect 23826 31955 24018 32059
rect 115 31937 364 31955
rect 50 31801 364 31937
rect 23648 31948 24018 31955
rect 23648 31902 23899 31948
rect 23945 31902 24018 31948
rect 23648 31801 24018 31902
rect 23826 30552 24018 30598
rect 23826 30506 23899 30552
rect 23945 30506 24018 30552
rect 50 30418 134 30437
rect 50 30278 69 30418
rect 115 30413 134 30418
rect 23826 30413 24018 30506
rect 115 30278 364 30413
rect 50 30259 364 30278
rect 23702 30388 24018 30413
rect 23702 30342 23899 30388
rect 23945 30342 24018 30388
rect 23702 30259 24018 30342
rect 361 29803 834 29858
rect 361 29757 414 29803
rect 460 29757 735 29803
rect 781 29757 834 29803
rect 361 29649 834 29757
rect 980 29803 1453 29858
rect 980 29757 1033 29803
rect 1079 29757 1354 29803
rect 1400 29757 1453 29803
rect 980 29649 1453 29757
rect 1599 29803 2072 29858
rect 1599 29757 1652 29803
rect 1698 29757 1973 29803
rect 2019 29757 2072 29803
rect 1599 29649 2072 29757
rect 2218 29803 2691 29858
rect 2218 29757 2271 29803
rect 2317 29757 2592 29803
rect 2638 29757 2691 29803
rect 2218 29649 2691 29757
rect 2837 29803 3310 29858
rect 2837 29757 2890 29803
rect 2936 29757 3211 29803
rect 3257 29757 3310 29803
rect 2837 29649 3310 29757
rect 3456 29803 3929 29858
rect 3456 29757 3509 29803
rect 3555 29757 3830 29803
rect 3876 29757 3929 29803
rect 3456 29649 3929 29757
rect 4075 29803 4548 29858
rect 4075 29757 4128 29803
rect 4174 29757 4449 29803
rect 4495 29757 4548 29803
rect 4075 29649 4548 29757
rect 4694 29803 5167 29858
rect 4694 29757 4747 29803
rect 4793 29757 5068 29803
rect 5114 29757 5167 29803
rect 4694 29649 5167 29757
rect 5313 29803 5786 29858
rect 5313 29757 5366 29803
rect 5412 29757 5687 29803
rect 5733 29757 5786 29803
rect 5313 29649 5786 29757
rect 5932 29803 6405 29858
rect 5932 29757 5985 29803
rect 6031 29757 6306 29803
rect 6352 29757 6405 29803
rect 5932 29649 6405 29757
rect 6551 29803 7024 29858
rect 6551 29757 6604 29803
rect 6650 29757 6925 29803
rect 6971 29757 7024 29803
rect 6551 29649 7024 29757
rect 7170 29803 7643 29858
rect 7170 29757 7223 29803
rect 7269 29757 7544 29803
rect 7590 29757 7643 29803
rect 7170 29649 7643 29757
rect 7789 29803 8262 29858
rect 7789 29757 7842 29803
rect 7888 29757 8163 29803
rect 8209 29757 8262 29803
rect 7789 29649 8262 29757
rect 8408 29803 8881 29858
rect 8408 29757 8461 29803
rect 8507 29757 8782 29803
rect 8828 29757 8881 29803
rect 8408 29649 8881 29757
rect 9027 29803 9500 29858
rect 9027 29757 9080 29803
rect 9126 29757 9401 29803
rect 9447 29757 9500 29803
rect 9027 29649 9500 29757
rect 9646 29803 10119 29858
rect 9646 29757 9699 29803
rect 9745 29757 10020 29803
rect 10066 29757 10119 29803
rect 9646 29649 10119 29757
rect 10265 29803 10738 29858
rect 10265 29757 10318 29803
rect 10364 29757 10639 29803
rect 10685 29757 10738 29803
rect 10265 29649 10738 29757
rect 10884 29803 11357 29858
rect 10884 29757 10937 29803
rect 10983 29757 11258 29803
rect 11304 29757 11357 29803
rect 10884 29649 11357 29757
rect 11503 29803 11976 29858
rect 11503 29757 11556 29803
rect 11602 29757 11877 29803
rect 11923 29757 11976 29803
rect 11503 29649 11976 29757
rect 12122 29803 12595 29858
rect 12122 29757 12175 29803
rect 12221 29757 12496 29803
rect 12542 29757 12595 29803
rect 12122 29649 12595 29757
rect 12741 29803 13214 29858
rect 12741 29757 12794 29803
rect 12840 29757 13115 29803
rect 13161 29757 13214 29803
rect 12741 29649 13214 29757
rect 13360 29803 13833 29858
rect 13360 29757 13413 29803
rect 13459 29757 13734 29803
rect 13780 29757 13833 29803
rect 13360 29649 13833 29757
rect 13979 29803 14452 29858
rect 13979 29757 14032 29803
rect 14078 29757 14353 29803
rect 14399 29757 14452 29803
rect 13979 29649 14452 29757
rect 14598 29803 15071 29858
rect 14598 29757 14651 29803
rect 14697 29757 14972 29803
rect 15018 29757 15071 29803
rect 14598 29649 15071 29757
rect 15217 29803 15690 29858
rect 15217 29757 15270 29803
rect 15316 29757 15591 29803
rect 15637 29757 15690 29803
rect 15217 29649 15690 29757
rect 15836 29803 16309 29858
rect 15836 29757 15889 29803
rect 15935 29757 16210 29803
rect 16256 29757 16309 29803
rect 15836 29649 16309 29757
rect 16455 29803 16928 29858
rect 16455 29757 16508 29803
rect 16554 29757 16829 29803
rect 16875 29757 16928 29803
rect 16455 29649 16928 29757
rect 17074 29803 17547 29858
rect 17074 29757 17127 29803
rect 17173 29757 17448 29803
rect 17494 29757 17547 29803
rect 17074 29649 17547 29757
rect 17693 29803 18166 29858
rect 17693 29757 17746 29803
rect 17792 29757 18067 29803
rect 18113 29757 18166 29803
rect 17693 29649 18166 29757
rect 18312 29803 18785 29858
rect 18312 29757 18365 29803
rect 18411 29757 18686 29803
rect 18732 29757 18785 29803
rect 18312 29649 18785 29757
rect 18931 29803 19404 29858
rect 18931 29757 18984 29803
rect 19030 29757 19305 29803
rect 19351 29757 19404 29803
rect 18931 29649 19404 29757
rect 19550 29803 20023 29858
rect 19550 29757 19603 29803
rect 19649 29757 19924 29803
rect 19970 29757 20023 29803
rect 19550 29649 20023 29757
rect 20169 29803 20642 29858
rect 20169 29757 20222 29803
rect 20268 29757 20543 29803
rect 20589 29757 20642 29803
rect 20169 29649 20642 29757
rect 20788 29803 21261 29858
rect 20788 29757 20841 29803
rect 20887 29757 21162 29803
rect 21208 29757 21261 29803
rect 20788 29649 21261 29757
rect 21407 29803 21880 29858
rect 21407 29757 21460 29803
rect 21506 29757 21781 29803
rect 21827 29757 21880 29803
rect 21407 29649 21880 29757
rect 22026 29803 22499 29858
rect 22026 29757 22079 29803
rect 22125 29757 22400 29803
rect 22446 29757 22499 29803
rect 22026 29649 22499 29757
rect 361 29112 834 29194
rect 980 29112 1453 29194
rect 1599 29112 2072 29194
rect 2218 29112 2691 29194
rect 2837 29112 3310 29194
rect 3456 29112 3929 29194
rect 4075 29112 4548 29194
rect 4694 29112 5167 29194
rect 5313 29112 5786 29194
rect 5932 29112 6405 29194
rect 6551 29112 7024 29194
rect 7170 29112 7643 29194
rect 7789 29112 8262 29194
rect 8408 29112 8881 29194
rect 9027 29112 9500 29194
rect 9646 29112 10119 29194
rect 10265 29112 10738 29194
rect 10884 29112 11357 29194
rect 11503 29112 11976 29194
rect 12122 29112 12595 29194
rect 12741 29112 13214 29194
rect 13360 29112 13833 29194
rect 13979 29112 14452 29194
rect 14598 29112 15071 29194
rect 15217 29112 15690 29194
rect 15836 29112 16309 29194
rect 16455 29112 16928 29194
rect 17074 29112 17547 29194
rect 17693 29112 18166 29194
rect 18312 29112 18785 29194
rect 18931 29112 19404 29194
rect 19550 29112 20023 29194
rect 20169 29112 20642 29194
rect 20788 29112 21261 29194
rect 21407 29112 21880 29194
rect 22026 29112 22499 29194
rect 23220 28632 23340 28705
rect 23444 28632 23564 28705
rect 23220 27857 23340 27950
rect 23444 27857 23564 27950
rect 23220 27115 23340 27175
rect 23444 27115 23564 27175
rect 23220 27093 23564 27115
rect 23220 27047 23328 27093
rect 23468 27047 23564 27093
rect 23220 27028 23564 27047
rect 23334 26956 23454 27028
rect 23334 25550 23454 25594
rect 23332 25369 23452 25413
rect 23332 23926 23452 24007
rect 23332 23880 23369 23926
rect 23415 23880 23452 23926
rect 23332 23861 23452 23880
rect 23332 23678 23452 23722
rect 23332 21674 23452 22316
rect 23332 20228 23452 20312
rect 23332 20182 23369 20228
rect 23415 20182 23452 20228
rect 23332 20163 23452 20182
rect 23332 19951 23452 19970
rect 23332 19905 23369 19951
rect 23415 19905 23452 19951
rect 23332 19819 23452 19905
rect 23332 18413 23452 18457
rect 23263 17984 23635 18003
rect 23263 17938 23426 17984
rect 23472 17938 23635 17984
rect 23263 17904 23635 17938
rect 23263 17844 23383 17904
rect 23515 17844 23635 17904
rect 23263 17360 23383 17547
rect 23515 17378 23635 17547
rect 23292 17329 23383 17360
rect 23516 17371 23635 17378
rect 23292 17256 23412 17329
rect 23516 17256 23636 17371
rect 23292 17069 23412 17142
rect 23516 17069 23636 17142
rect 23243 15171 23363 15215
rect 23467 15171 23587 15215
rect 23243 14409 23363 14469
rect 23467 14409 23587 14469
rect 23243 14393 23587 14409
rect 23243 14347 23876 14393
rect 23243 14301 23598 14347
rect 23644 14301 23756 14347
rect 23802 14301 23876 14347
rect 23243 14255 23876 14301
rect 23243 14246 23587 14255
rect 23243 14165 23363 14246
rect 23467 14165 23587 14246
rect 23243 13806 23363 13889
rect 23467 13806 23587 13889
rect 23247 12504 23367 12548
rect 23471 12504 23591 12548
rect 23247 10741 23367 10804
rect 23471 10741 23591 10804
rect 23247 10732 23591 10741
rect 22940 10686 23591 10732
rect 22940 10640 23014 10686
rect 23060 10640 23172 10686
rect 23218 10640 23591 10686
rect 22940 10594 23591 10640
rect 23247 10583 23591 10594
rect 23247 10523 23367 10583
rect 23471 10523 23591 10583
rect 23247 8351 23367 8395
rect 23471 8351 23591 8395
<< polycontact >>
rect 69 89396 115 89536
rect 23899 89426 23945 89472
rect 23899 89262 23945 89308
rect 69 87737 115 87877
rect 23899 87866 23945 87912
rect 23899 87702 23945 87748
rect 69 85937 115 86077
rect 23899 86066 23945 86112
rect 23899 85902 23945 85948
rect 69 84137 115 84277
rect 23899 84266 23945 84312
rect 23899 84102 23945 84148
rect 69 82337 115 82477
rect 23899 82466 23945 82512
rect 23899 82302 23945 82348
rect 69 80537 115 80677
rect 23899 80666 23945 80712
rect 23899 80502 23945 80548
rect 69 78737 115 78877
rect 23899 78866 23945 78912
rect 23899 78702 23945 78748
rect 69 76937 115 77077
rect 23899 77066 23945 77112
rect 23899 76902 23945 76948
rect 69 75137 115 75277
rect 23899 75266 23945 75312
rect 23899 75102 23945 75148
rect 69 73337 115 73477
rect 23899 73466 23945 73512
rect 23899 73302 23945 73348
rect 69 71537 115 71677
rect 23899 71666 23945 71712
rect 23899 71502 23945 71548
rect 69 69737 115 69877
rect 23899 69866 23945 69912
rect 23899 69702 23945 69748
rect 69 67937 115 68077
rect 23899 68066 23945 68112
rect 23899 67902 23945 67948
rect 69 66137 115 66277
rect 23899 66266 23945 66312
rect 23899 66102 23945 66148
rect 69 64337 115 64477
rect 23899 64466 23945 64512
rect 23899 64302 23945 64348
rect 69 62537 115 62677
rect 23899 62666 23945 62712
rect 23899 62502 23945 62548
rect 69 60737 115 60877
rect 23899 60866 23945 60912
rect 23899 60702 23945 60748
rect 69 58937 115 59077
rect 23899 59066 23945 59112
rect 23899 58902 23945 58948
rect 69 57137 115 57277
rect 23899 57266 23945 57312
rect 23899 57102 23945 57148
rect 69 55337 115 55477
rect 23899 55466 23945 55512
rect 23899 55302 23945 55348
rect 69 53537 115 53677
rect 23899 53666 23945 53712
rect 23899 53502 23945 53548
rect 69 51737 115 51877
rect 23899 51866 23945 51912
rect 23899 51702 23945 51748
rect 69 49937 115 50077
rect 23899 50066 23945 50112
rect 23899 49902 23945 49948
rect 69 48137 115 48277
rect 23899 48266 23945 48312
rect 23899 48102 23945 48148
rect 69 46337 115 46477
rect 23899 46466 23945 46512
rect 23899 46302 23945 46348
rect 69 44537 115 44677
rect 23899 44666 23945 44712
rect 23899 44502 23945 44548
rect 69 42737 115 42877
rect 23899 42866 23945 42912
rect 23899 42702 23945 42748
rect 69 40937 115 41077
rect 23899 41066 23945 41112
rect 23899 40902 23945 40948
rect 69 39137 115 39277
rect 23899 39266 23945 39312
rect 23899 39102 23945 39148
rect 69 37337 115 37477
rect 23899 37466 23945 37512
rect 23899 37302 23945 37348
rect 69 35537 115 35677
rect 23899 35666 23945 35712
rect 23899 35502 23945 35548
rect 69 33737 115 33877
rect 23899 33866 23945 33912
rect 23899 33702 23945 33748
rect 69 31937 115 32077
rect 23899 32066 23945 32112
rect 23899 31902 23945 31948
rect 23899 30506 23945 30552
rect 69 30278 115 30418
rect 23899 30342 23945 30388
rect 414 29757 460 29803
rect 735 29757 781 29803
rect 1033 29757 1079 29803
rect 1354 29757 1400 29803
rect 1652 29757 1698 29803
rect 1973 29757 2019 29803
rect 2271 29757 2317 29803
rect 2592 29757 2638 29803
rect 2890 29757 2936 29803
rect 3211 29757 3257 29803
rect 3509 29757 3555 29803
rect 3830 29757 3876 29803
rect 4128 29757 4174 29803
rect 4449 29757 4495 29803
rect 4747 29757 4793 29803
rect 5068 29757 5114 29803
rect 5366 29757 5412 29803
rect 5687 29757 5733 29803
rect 5985 29757 6031 29803
rect 6306 29757 6352 29803
rect 6604 29757 6650 29803
rect 6925 29757 6971 29803
rect 7223 29757 7269 29803
rect 7544 29757 7590 29803
rect 7842 29757 7888 29803
rect 8163 29757 8209 29803
rect 8461 29757 8507 29803
rect 8782 29757 8828 29803
rect 9080 29757 9126 29803
rect 9401 29757 9447 29803
rect 9699 29757 9745 29803
rect 10020 29757 10066 29803
rect 10318 29757 10364 29803
rect 10639 29757 10685 29803
rect 10937 29757 10983 29803
rect 11258 29757 11304 29803
rect 11556 29757 11602 29803
rect 11877 29757 11923 29803
rect 12175 29757 12221 29803
rect 12496 29757 12542 29803
rect 12794 29757 12840 29803
rect 13115 29757 13161 29803
rect 13413 29757 13459 29803
rect 13734 29757 13780 29803
rect 14032 29757 14078 29803
rect 14353 29757 14399 29803
rect 14651 29757 14697 29803
rect 14972 29757 15018 29803
rect 15270 29757 15316 29803
rect 15591 29757 15637 29803
rect 15889 29757 15935 29803
rect 16210 29757 16256 29803
rect 16508 29757 16554 29803
rect 16829 29757 16875 29803
rect 17127 29757 17173 29803
rect 17448 29757 17494 29803
rect 17746 29757 17792 29803
rect 18067 29757 18113 29803
rect 18365 29757 18411 29803
rect 18686 29757 18732 29803
rect 18984 29757 19030 29803
rect 19305 29757 19351 29803
rect 19603 29757 19649 29803
rect 19924 29757 19970 29803
rect 20222 29757 20268 29803
rect 20543 29757 20589 29803
rect 20841 29757 20887 29803
rect 21162 29757 21208 29803
rect 21460 29757 21506 29803
rect 21781 29757 21827 29803
rect 22079 29757 22125 29803
rect 22400 29757 22446 29803
rect 23328 27047 23468 27093
rect 23369 23880 23415 23926
rect 23369 20182 23415 20228
rect 23369 19905 23415 19951
rect 23426 17938 23472 17984
rect 23598 14301 23644 14347
rect 23756 14301 23802 14347
rect 23014 10640 23060 10686
rect 23172 10640 23218 10686
<< metal1 >>
rect 54 89536 130 89547
rect 54 89535 69 89536
rect 115 89535 130 89536
rect 54 89275 66 89535
rect 118 89275 130 89535
rect 54 89263 130 89275
rect 23858 89477 23982 89517
rect 23858 89425 23894 89477
rect 23946 89425 23982 89477
rect 23858 89308 23982 89425
rect 23858 89262 23899 89308
rect 23945 89262 23982 89308
rect 23858 89259 23982 89262
rect 23858 89207 23894 89259
rect 23946 89207 23982 89259
rect 23858 89167 23982 89207
rect 54 87936 130 87948
rect 54 87676 66 87936
rect 118 87676 130 87936
rect 54 87664 130 87676
rect 23858 87940 23982 87980
rect 23858 87888 23894 87940
rect 23946 87888 23982 87940
rect 23858 87866 23899 87888
rect 23945 87866 23982 87888
rect 23858 87748 23982 87866
rect 23858 87722 23899 87748
rect 23945 87722 23982 87748
rect 23858 87670 23894 87722
rect 23946 87670 23982 87722
rect 23858 87630 23982 87670
rect 54 86137 130 86149
rect 54 85877 66 86137
rect 118 85877 130 86137
rect 54 85865 130 85877
rect 23858 86140 23982 86180
rect 23858 86088 23894 86140
rect 23946 86088 23982 86140
rect 23858 86066 23899 86088
rect 23945 86066 23982 86088
rect 23858 85948 23982 86066
rect 23858 85922 23899 85948
rect 23945 85922 23982 85948
rect 23858 85870 23894 85922
rect 23946 85870 23982 85922
rect 23858 85830 23982 85870
rect 54 84337 130 84349
rect 54 84077 66 84337
rect 118 84077 130 84337
rect 54 84065 130 84077
rect 23858 84340 23982 84380
rect 23858 84288 23894 84340
rect 23946 84288 23982 84340
rect 23858 84266 23899 84288
rect 23945 84266 23982 84288
rect 23858 84148 23982 84266
rect 23858 84122 23899 84148
rect 23945 84122 23982 84148
rect 23858 84070 23894 84122
rect 23946 84070 23982 84122
rect 23858 84030 23982 84070
rect 54 82537 130 82549
rect 54 82277 66 82537
rect 118 82277 130 82537
rect 54 82265 130 82277
rect 23858 82540 23982 82580
rect 23858 82488 23894 82540
rect 23946 82488 23982 82540
rect 23858 82466 23899 82488
rect 23945 82466 23982 82488
rect 23858 82348 23982 82466
rect 23858 82322 23899 82348
rect 23945 82322 23982 82348
rect 23858 82270 23894 82322
rect 23946 82270 23982 82322
rect 23858 82230 23982 82270
rect 54 80736 130 80748
rect 54 80476 66 80736
rect 118 80476 130 80736
rect 54 80464 130 80476
rect 23858 80740 23982 80780
rect 23858 80688 23894 80740
rect 23946 80707 23982 80740
rect 23946 80688 24405 80707
rect 23858 80666 23899 80688
rect 23945 80666 24405 80688
rect 23858 80548 24405 80666
rect 23858 80522 23899 80548
rect 23945 80522 24405 80548
rect 23858 80470 23894 80522
rect 23946 80507 24405 80522
rect 23946 80470 23982 80507
rect 23858 80430 23982 80470
rect 54 78937 130 78949
rect 54 78677 66 78937
rect 118 78677 130 78937
rect 54 78665 130 78677
rect 23858 78940 23982 78980
rect 23858 78888 23894 78940
rect 23946 78888 23982 78940
rect 23858 78866 23899 78888
rect 23945 78866 23982 78888
rect 23858 78748 23982 78866
rect 23858 78722 23899 78748
rect 23945 78722 23982 78748
rect 23858 78670 23894 78722
rect 23946 78670 23982 78722
rect 23858 78630 23982 78670
rect 54 77138 130 77150
rect 54 76878 66 77138
rect 118 76878 130 77138
rect 54 76866 130 76878
rect 23858 77140 23982 77180
rect 23858 77088 23894 77140
rect 23946 77088 23982 77140
rect 23858 77066 23899 77088
rect 23945 77066 23982 77088
rect 23858 76948 23982 77066
rect 23858 76922 23899 76948
rect 23945 76922 23982 76948
rect 23858 76870 23894 76922
rect 23946 76870 23982 76922
rect 23858 76830 23982 76870
rect 54 75337 130 75349
rect 54 75077 66 75337
rect 118 75077 130 75337
rect 54 75065 130 75077
rect 23858 75340 23982 75380
rect 23858 75288 23894 75340
rect 23946 75288 23982 75340
rect 23858 75266 23899 75288
rect 23945 75266 23982 75288
rect 23858 75148 23982 75266
rect 23858 75122 23899 75148
rect 23945 75122 23982 75148
rect 23858 75070 23894 75122
rect 23946 75070 23982 75122
rect 23858 75030 23982 75070
rect 54 73537 130 73549
rect 54 73277 66 73537
rect 118 73277 130 73537
rect 54 73265 130 73277
rect 23858 73540 23982 73580
rect 23858 73488 23894 73540
rect 23946 73488 23982 73540
rect 23858 73466 23899 73488
rect 23945 73466 23982 73488
rect 23858 73348 23982 73466
rect 23858 73322 23899 73348
rect 23945 73322 23982 73348
rect 23858 73270 23894 73322
rect 23946 73270 23982 73322
rect 23858 73230 23982 73270
rect 54 71737 130 71749
rect 54 71477 66 71737
rect 118 71477 130 71737
rect 54 71465 130 71477
rect 23858 71740 23982 71780
rect 23858 71688 23894 71740
rect 23946 71688 23982 71740
rect 23858 71666 23899 71688
rect 23945 71666 23982 71688
rect 23858 71548 23982 71666
rect 23858 71522 23899 71548
rect 23945 71522 23982 71548
rect 23858 71470 23894 71522
rect 23946 71470 23982 71522
rect 23858 71430 23982 71470
rect 54 69937 130 69949
rect 54 69677 66 69937
rect 118 69677 130 69937
rect 54 69665 130 69677
rect 23858 69940 23982 69980
rect 23858 69888 23894 69940
rect 23946 69888 23982 69940
rect 23858 69866 23899 69888
rect 23945 69866 23982 69888
rect 23858 69748 23982 69866
rect 23858 69722 23899 69748
rect 23945 69722 23982 69748
rect 23858 69670 23894 69722
rect 23946 69670 23982 69722
rect 23858 69630 23982 69670
rect 54 68137 130 68149
rect 54 67877 66 68137
rect 118 67877 130 68137
rect 54 67865 130 67877
rect 23858 68140 23982 68180
rect 23858 68088 23894 68140
rect 23946 68088 23982 68140
rect 23858 68066 23899 68088
rect 23945 68066 23982 68088
rect 23858 67948 23982 68066
rect 23858 67922 23899 67948
rect 23945 67922 23982 67948
rect 23858 67870 23894 67922
rect 23946 67870 23982 67922
rect 23858 67830 23982 67870
rect 54 66337 130 66349
rect 54 66077 66 66337
rect 118 66077 130 66337
rect 54 66065 130 66077
rect 23858 66340 23982 66380
rect 23858 66288 23894 66340
rect 23946 66288 23982 66340
rect 23858 66266 23899 66288
rect 23945 66266 23982 66288
rect 23858 66148 23982 66266
rect 23858 66122 23899 66148
rect 23945 66122 23982 66148
rect 23858 66070 23894 66122
rect 23946 66070 23982 66122
rect 23858 66030 23982 66070
rect 54 64537 130 64549
rect 54 64277 66 64537
rect 118 64277 130 64537
rect 54 64265 130 64277
rect 23858 64540 23982 64580
rect 23858 64488 23894 64540
rect 23946 64488 23982 64540
rect 23858 64466 23899 64488
rect 23945 64466 23982 64488
rect 23858 64348 23982 64466
rect 23858 64322 23899 64348
rect 23945 64322 23982 64348
rect 23858 64270 23894 64322
rect 23946 64270 23982 64322
rect 23858 64230 23982 64270
rect 54 62737 130 62749
rect 54 62477 66 62737
rect 118 62477 130 62737
rect 54 62465 130 62477
rect 23858 62740 23982 62780
rect 23858 62688 23894 62740
rect 23946 62688 23982 62740
rect 23858 62666 23899 62688
rect 23945 62666 23982 62688
rect 23858 62548 23982 62666
rect 23858 62522 23899 62548
rect 23945 62522 23982 62548
rect 23858 62470 23894 62522
rect 23946 62470 23982 62522
rect 23858 62430 23982 62470
rect 54 60937 130 60949
rect 54 60677 66 60937
rect 118 60677 130 60937
rect 54 60665 130 60677
rect 23858 60940 23982 60980
rect 23858 60888 23894 60940
rect 23946 60888 23982 60940
rect 23858 60866 23899 60888
rect 23945 60866 23982 60888
rect 23858 60748 23982 60866
rect 23858 60722 23899 60748
rect 23945 60722 23982 60748
rect 23858 60670 23894 60722
rect 23946 60670 23982 60722
rect 23858 60630 23982 60670
rect 54 59137 130 59149
rect 54 58877 66 59137
rect 118 58877 130 59137
rect 54 58865 130 58877
rect 23858 59140 23982 59180
rect 23858 59088 23894 59140
rect 23946 59088 23982 59140
rect 23858 59066 23899 59088
rect 23945 59066 23982 59088
rect 23858 58948 23982 59066
rect 23858 58922 23899 58948
rect 23945 58922 23982 58948
rect 23858 58870 23894 58922
rect 23946 58870 23982 58922
rect 23858 58830 23982 58870
rect 54 57337 130 57349
rect 54 57077 66 57337
rect 118 57077 130 57337
rect 54 57065 130 57077
rect 23858 57340 23982 57380
rect 23858 57288 23894 57340
rect 23946 57288 23982 57340
rect 23858 57266 23899 57288
rect 23945 57266 23982 57288
rect 23858 57148 23982 57266
rect 23858 57122 23899 57148
rect 23945 57122 23982 57148
rect 23858 57070 23894 57122
rect 23946 57070 23982 57122
rect 23858 57030 23982 57070
rect 54 55537 130 55549
rect 54 55277 66 55537
rect 118 55277 130 55537
rect 54 55265 130 55277
rect 23858 55544 23982 55584
rect 23858 55492 23894 55544
rect 23946 55492 23982 55544
rect 23858 55466 23899 55492
rect 23945 55466 23982 55492
rect 23858 55348 23982 55466
rect 23858 55326 23899 55348
rect 23945 55326 23982 55348
rect 23858 55274 23894 55326
rect 23946 55274 23982 55326
rect 23858 55234 23982 55274
rect 50 53737 126 53749
rect 50 53477 62 53737
rect 114 53677 126 53737
rect 115 53537 126 53677
rect 114 53477 126 53537
rect 50 53465 126 53477
rect 23858 53740 23982 53780
rect 23858 53688 23894 53740
rect 23946 53688 23982 53740
rect 23858 53666 23899 53688
rect 23945 53666 23982 53688
rect 23858 53548 23982 53666
rect 23858 53522 23899 53548
rect 23945 53522 23982 53548
rect 23858 53470 23894 53522
rect 23946 53470 23982 53522
rect 23858 53430 23982 53470
rect 54 51937 130 51949
rect 54 51677 66 51937
rect 118 51677 130 51937
rect 54 51665 130 51677
rect 23858 51944 23982 51984
rect 23858 51892 23894 51944
rect 23946 51892 23982 51944
rect 23858 51866 23899 51892
rect 23945 51866 23982 51892
rect 23858 51748 23982 51866
rect 23858 51726 23899 51748
rect 23945 51726 23982 51748
rect 23858 51674 23894 51726
rect 23946 51674 23982 51726
rect 23858 51634 23982 51674
rect 54 50137 130 50149
rect 54 49877 66 50137
rect 118 49877 130 50137
rect 54 49865 130 49877
rect 23858 50140 23982 50180
rect 23858 50088 23894 50140
rect 23946 50088 23982 50140
rect 23858 50066 23899 50088
rect 23945 50066 23982 50088
rect 23858 49948 23982 50066
rect 23858 49922 23899 49948
rect 23945 49922 23982 49948
rect 23858 49870 23894 49922
rect 23946 49870 23982 49922
rect 23858 49830 23982 49870
rect 54 48337 130 48349
rect 54 48077 66 48337
rect 118 48077 130 48337
rect 54 48065 130 48077
rect 23858 48344 23982 48384
rect 23858 48292 23894 48344
rect 23946 48292 23982 48344
rect 23858 48266 23899 48292
rect 23945 48266 23982 48292
rect 23858 48148 23982 48266
rect 23858 48126 23899 48148
rect 23945 48126 23982 48148
rect 23858 48074 23894 48126
rect 23946 48074 23982 48126
rect 23858 48034 23982 48074
rect 54 46537 130 46549
rect 54 46277 66 46537
rect 118 46277 130 46537
rect 54 46265 130 46277
rect 23858 46540 23982 46580
rect 23858 46488 23894 46540
rect 23946 46488 23982 46540
rect 23858 46466 23899 46488
rect 23945 46466 23982 46488
rect 23858 46348 23982 46466
rect 23858 46322 23899 46348
rect 23945 46322 23982 46348
rect 23858 46270 23894 46322
rect 23946 46270 23982 46322
rect 23858 46230 23982 46270
rect 54 44737 130 44749
rect 54 44477 66 44737
rect 118 44477 130 44737
rect 54 44465 130 44477
rect 23858 44744 23982 44784
rect 23858 44692 23894 44744
rect 23946 44692 23982 44744
rect 23858 44666 23899 44692
rect 23945 44666 23982 44692
rect 23858 44548 23982 44666
rect 23858 44526 23899 44548
rect 23945 44526 23982 44548
rect 23858 44474 23894 44526
rect 23946 44474 23982 44526
rect 23858 44434 23982 44474
rect 54 42937 130 42949
rect 54 42677 66 42937
rect 118 42677 130 42937
rect 54 42665 130 42677
rect 23858 42940 23982 42980
rect 23858 42888 23894 42940
rect 23946 42888 23982 42940
rect 23858 42866 23899 42888
rect 23945 42866 23982 42888
rect 23858 42748 23982 42866
rect 23858 42722 23899 42748
rect 23945 42722 23982 42748
rect 23858 42670 23894 42722
rect 23946 42670 23982 42722
rect 23858 42630 23982 42670
rect 54 41137 130 41149
rect 54 40877 66 41137
rect 118 40877 130 41137
rect 54 40865 130 40877
rect 23858 41144 23982 41184
rect 23858 41092 23894 41144
rect 23946 41092 23982 41144
rect 23858 41066 23899 41092
rect 23945 41066 23982 41092
rect 23858 40948 23982 41066
rect 23858 40926 23899 40948
rect 23945 40926 23982 40948
rect 23858 40874 23894 40926
rect 23946 40874 23982 40926
rect 23858 40834 23982 40874
rect 54 39337 130 39349
rect 54 39077 66 39337
rect 118 39077 130 39337
rect 54 39065 130 39077
rect 23858 39340 23982 39380
rect 23858 39288 23894 39340
rect 23946 39288 23982 39340
rect 23858 39266 23899 39288
rect 23945 39266 23982 39288
rect 23858 39148 23982 39266
rect 23858 39122 23899 39148
rect 23945 39122 23982 39148
rect 23858 39070 23894 39122
rect 23946 39070 23982 39122
rect 23858 39030 23982 39070
rect 54 37537 130 37549
rect 54 37277 66 37537
rect 118 37277 130 37537
rect 54 37265 130 37277
rect 23858 37544 23982 37584
rect 23858 37492 23894 37544
rect 23946 37492 23982 37544
rect 23858 37466 23899 37492
rect 23945 37466 23982 37492
rect 23858 37348 23982 37466
rect 23858 37326 23899 37348
rect 23945 37326 23982 37348
rect 23858 37274 23894 37326
rect 23946 37274 23982 37326
rect 23858 37234 23982 37274
rect 54 35737 130 35749
rect 54 35477 66 35737
rect 118 35477 130 35737
rect 54 35465 130 35477
rect 23858 35740 23982 35780
rect 23858 35688 23894 35740
rect 23946 35688 23982 35740
rect 23858 35666 23899 35688
rect 23945 35666 23982 35688
rect 23858 35548 23982 35666
rect 23858 35522 23899 35548
rect 23945 35522 23982 35548
rect 23858 35470 23894 35522
rect 23946 35470 23982 35522
rect 23858 35430 23982 35470
rect 54 33937 130 33949
rect 54 33677 66 33937
rect 118 33677 130 33937
rect 54 33665 130 33677
rect 23858 33944 23982 33984
rect 23858 33892 23894 33944
rect 23946 33892 23982 33944
rect 23858 33866 23899 33892
rect 23945 33866 23982 33892
rect 23858 33748 23982 33866
rect 23858 33726 23899 33748
rect 23945 33726 23982 33748
rect 23858 33674 23894 33726
rect 23946 33674 23982 33726
rect 23858 33634 23982 33674
rect 54 32137 130 32149
rect 54 31877 66 32137
rect 118 31877 130 32137
rect 54 31865 130 31877
rect 23858 32140 23982 32180
rect 23858 32088 23894 32140
rect 23946 32088 23982 32140
rect 23858 32066 23899 32088
rect 23945 32066 23982 32088
rect 23858 31948 23982 32066
rect 23858 31922 23899 31948
rect 23945 31922 23982 31948
rect 23858 31870 23894 31922
rect 23946 31870 23982 31922
rect 23858 31830 23982 31870
rect 23858 30607 23982 30647
rect 23858 30555 23894 30607
rect 23946 30555 23982 30607
rect 23858 30552 23982 30555
rect 23858 30506 23899 30552
rect 23945 30506 23982 30552
rect 52 30418 128 30487
rect 52 30278 69 30418
rect 115 30278 128 30418
rect 23858 30389 23982 30506
rect 23858 30337 23894 30389
rect 23946 30337 23982 30389
rect 23858 30297 23982 30337
rect 52 29890 128 30278
rect 1125 29890 1289 30167
rect 6525 29890 6689 30167
rect 11925 29890 12089 30167
rect 17325 29890 17489 30167
rect 22725 29890 22889 30167
rect 52 29818 24835 29890
rect 52 29803 948 29818
rect 1104 29803 11742 29818
rect 11898 29803 22869 29818
rect 52 29757 414 29803
rect 460 29757 735 29803
rect 781 29766 948 29803
rect 1104 29766 1354 29803
rect 781 29757 1033 29766
rect 1079 29757 1354 29766
rect 1400 29757 1652 29803
rect 1698 29757 1973 29803
rect 2019 29757 2271 29803
rect 2317 29757 2592 29803
rect 2638 29757 2890 29803
rect 2936 29757 3211 29803
rect 3257 29757 3509 29803
rect 3555 29757 3830 29803
rect 3876 29757 4128 29803
rect 4174 29757 4449 29803
rect 4495 29757 4747 29803
rect 4793 29757 5068 29803
rect 5114 29757 5366 29803
rect 5412 29757 5687 29803
rect 5733 29757 5985 29803
rect 6031 29757 6306 29803
rect 6352 29757 6604 29803
rect 6650 29757 6925 29803
rect 6971 29757 7223 29803
rect 7269 29757 7544 29803
rect 7590 29757 7842 29803
rect 7888 29757 8163 29803
rect 8209 29757 8461 29803
rect 8507 29757 8782 29803
rect 8828 29757 9080 29803
rect 9126 29757 9401 29803
rect 9447 29757 9699 29803
rect 9745 29757 10020 29803
rect 10066 29757 10318 29803
rect 10364 29757 10639 29803
rect 10685 29757 10937 29803
rect 10983 29757 11258 29803
rect 11304 29757 11556 29803
rect 11602 29766 11742 29803
rect 11602 29757 11877 29766
rect 11923 29757 12175 29803
rect 12221 29757 12496 29803
rect 12542 29757 12794 29803
rect 12840 29757 13115 29803
rect 13161 29757 13413 29803
rect 13459 29757 13734 29803
rect 13780 29757 14032 29803
rect 14078 29757 14353 29803
rect 14399 29757 14651 29803
rect 14697 29757 14972 29803
rect 15018 29757 15270 29803
rect 15316 29757 15591 29803
rect 15637 29757 15889 29803
rect 15935 29757 16210 29803
rect 16256 29757 16508 29803
rect 16554 29757 16829 29803
rect 16875 29757 17127 29803
rect 17173 29757 17448 29803
rect 17494 29757 17746 29803
rect 17792 29757 18067 29803
rect 18113 29757 18365 29803
rect 18411 29757 18686 29803
rect 18732 29757 18984 29803
rect 19030 29757 19305 29803
rect 19351 29757 19603 29803
rect 19649 29757 19924 29803
rect 19970 29757 20222 29803
rect 20268 29757 20543 29803
rect 20589 29757 20841 29803
rect 20887 29757 21162 29803
rect 21208 29757 21460 29803
rect 21506 29757 21781 29803
rect 21827 29757 22079 29803
rect 22125 29757 22400 29803
rect 22446 29766 22869 29803
rect 23025 29766 24835 29818
rect 22446 29757 24835 29766
rect 52 29720 24835 29757
rect 230 29604 346 29640
rect 230 29558 265 29604
rect 311 29558 346 29604
rect 230 29286 346 29558
rect 230 29240 265 29286
rect 311 29240 346 29286
rect 230 28890 346 29240
rect 849 29604 965 29640
rect 849 29558 884 29604
rect 930 29558 965 29604
rect 849 29286 965 29558
rect 849 29240 884 29286
rect 930 29240 965 29286
rect 849 28890 965 29240
rect 1468 29604 1584 29640
rect 1468 29558 1503 29604
rect 1549 29558 1584 29604
rect 1468 29286 1584 29558
rect 1468 29240 1503 29286
rect 1549 29240 1584 29286
rect 1468 28890 1584 29240
rect 2087 29604 2203 29640
rect 2087 29558 2122 29604
rect 2168 29558 2203 29604
rect 2087 29286 2203 29558
rect 2087 29240 2122 29286
rect 2168 29240 2203 29286
rect 2087 28890 2203 29240
rect 2706 29604 2822 29640
rect 2706 29558 2741 29604
rect 2787 29558 2822 29604
rect 2706 29286 2822 29558
rect 2706 29240 2741 29286
rect 2787 29240 2822 29286
rect 2706 28890 2822 29240
rect 3325 29604 3441 29640
rect 3325 29558 3360 29604
rect 3406 29558 3441 29604
rect 3325 29286 3441 29558
rect 3325 29240 3360 29286
rect 3406 29240 3441 29286
rect 3325 28890 3441 29240
rect 3944 29604 4060 29640
rect 3944 29558 3979 29604
rect 4025 29558 4060 29604
rect 3944 29286 4060 29558
rect 3944 29240 3979 29286
rect 4025 29240 4060 29286
rect 3944 28890 4060 29240
rect 4563 29604 4679 29640
rect 4563 29558 4598 29604
rect 4644 29558 4679 29604
rect 4563 29286 4679 29558
rect 4563 29240 4598 29286
rect 4644 29240 4679 29286
rect 4563 28890 4679 29240
rect 5182 29604 5298 29640
rect 5182 29558 5217 29604
rect 5263 29558 5298 29604
rect 5182 29286 5298 29558
rect 5182 29240 5217 29286
rect 5263 29240 5298 29286
rect 5182 28890 5298 29240
rect 5801 29604 5917 29640
rect 5801 29558 5836 29604
rect 5882 29558 5917 29604
rect 5801 29286 5917 29558
rect 5801 29240 5836 29286
rect 5882 29240 5917 29286
rect 5801 28890 5917 29240
rect 6420 29604 6536 29640
rect 6420 29558 6455 29604
rect 6501 29558 6536 29604
rect 6420 29286 6536 29558
rect 6420 29240 6455 29286
rect 6501 29240 6536 29286
rect 6420 28890 6536 29240
rect 7039 29604 7155 29640
rect 7039 29558 7074 29604
rect 7120 29558 7155 29604
rect 7039 29286 7155 29558
rect 7039 29240 7074 29286
rect 7120 29240 7155 29286
rect 7039 28890 7155 29240
rect 7658 29604 7774 29640
rect 7658 29558 7693 29604
rect 7739 29558 7774 29604
rect 7658 29286 7774 29558
rect 7658 29240 7693 29286
rect 7739 29240 7774 29286
rect 7658 28890 7774 29240
rect 8277 29604 8393 29640
rect 8277 29558 8312 29604
rect 8358 29558 8393 29604
rect 8277 29286 8393 29558
rect 8277 29240 8312 29286
rect 8358 29240 8393 29286
rect 8277 28890 8393 29240
rect 8896 29604 9012 29640
rect 8896 29558 8931 29604
rect 8977 29558 9012 29604
rect 8896 29286 9012 29558
rect 8896 29240 8931 29286
rect 8977 29240 9012 29286
rect 8896 28890 9012 29240
rect 9515 29604 9631 29640
rect 9515 29558 9550 29604
rect 9596 29558 9631 29604
rect 9515 29286 9631 29558
rect 9515 29240 9550 29286
rect 9596 29240 9631 29286
rect 9515 28890 9631 29240
rect 10134 29604 10250 29640
rect 10134 29558 10169 29604
rect 10215 29558 10250 29604
rect 10134 29286 10250 29558
rect 10134 29240 10169 29286
rect 10215 29240 10250 29286
rect 10134 28890 10250 29240
rect 10753 29604 10869 29640
rect 10753 29558 10788 29604
rect 10834 29558 10869 29604
rect 10753 29286 10869 29558
rect 10753 29240 10788 29286
rect 10834 29240 10869 29286
rect 10753 28890 10869 29240
rect 11372 29604 11488 29640
rect 11372 29558 11407 29604
rect 11453 29558 11488 29604
rect 11372 29286 11488 29558
rect 11372 29240 11407 29286
rect 11453 29240 11488 29286
rect 11372 28890 11488 29240
rect 11991 29604 12107 29640
rect 11991 29558 12026 29604
rect 12072 29558 12107 29604
rect 11991 29286 12107 29558
rect 11991 29240 12026 29286
rect 12072 29240 12107 29286
rect 11991 28890 12107 29240
rect 12610 29604 12726 29640
rect 12610 29558 12645 29604
rect 12691 29558 12726 29604
rect 12610 29286 12726 29558
rect 12610 29240 12645 29286
rect 12691 29240 12726 29286
rect 12610 28890 12726 29240
rect 13229 29604 13345 29640
rect 13229 29558 13264 29604
rect 13310 29558 13345 29604
rect 13229 29286 13345 29558
rect 13229 29240 13264 29286
rect 13310 29240 13345 29286
rect 13229 28890 13345 29240
rect 13848 29604 13964 29640
rect 13848 29558 13883 29604
rect 13929 29558 13964 29604
rect 13848 29286 13964 29558
rect 13848 29240 13883 29286
rect 13929 29240 13964 29286
rect 13848 28890 13964 29240
rect 14467 29604 14583 29640
rect 14467 29558 14502 29604
rect 14548 29558 14583 29604
rect 14467 29286 14583 29558
rect 14467 29240 14502 29286
rect 14548 29240 14583 29286
rect 14467 28890 14583 29240
rect 15086 29604 15202 29640
rect 15086 29558 15121 29604
rect 15167 29558 15202 29604
rect 15086 29286 15202 29558
rect 15086 29240 15121 29286
rect 15167 29240 15202 29286
rect 15086 28890 15202 29240
rect 15705 29604 15821 29640
rect 15705 29558 15740 29604
rect 15786 29558 15821 29604
rect 15705 29286 15821 29558
rect 15705 29240 15740 29286
rect 15786 29240 15821 29286
rect 15705 28890 15821 29240
rect 16324 29604 16440 29640
rect 16324 29558 16359 29604
rect 16405 29558 16440 29604
rect 16324 29286 16440 29558
rect 16324 29240 16359 29286
rect 16405 29240 16440 29286
rect 16324 28890 16440 29240
rect 16943 29604 17059 29640
rect 16943 29558 16978 29604
rect 17024 29558 17059 29604
rect 16943 29286 17059 29558
rect 16943 29240 16978 29286
rect 17024 29240 17059 29286
rect 16943 28890 17059 29240
rect 17562 29604 17678 29640
rect 17562 29558 17597 29604
rect 17643 29558 17678 29604
rect 17562 29286 17678 29558
rect 17562 29240 17597 29286
rect 17643 29240 17678 29286
rect 17562 28890 17678 29240
rect 18181 29604 18297 29640
rect 18181 29558 18216 29604
rect 18262 29558 18297 29604
rect 18181 29286 18297 29558
rect 18181 29240 18216 29286
rect 18262 29240 18297 29286
rect 18181 28890 18297 29240
rect 18800 29604 18916 29640
rect 18800 29558 18835 29604
rect 18881 29558 18916 29604
rect 18800 29286 18916 29558
rect 18800 29240 18835 29286
rect 18881 29240 18916 29286
rect 18800 28890 18916 29240
rect 19419 29604 19535 29640
rect 19419 29558 19454 29604
rect 19500 29558 19535 29604
rect 19419 29286 19535 29558
rect 19419 29240 19454 29286
rect 19500 29240 19535 29286
rect 19419 28890 19535 29240
rect 20038 29604 20154 29640
rect 20038 29558 20073 29604
rect 20119 29558 20154 29604
rect 20038 29286 20154 29558
rect 20038 29240 20073 29286
rect 20119 29240 20154 29286
rect 20038 28890 20154 29240
rect 20657 29604 20773 29640
rect 20657 29558 20692 29604
rect 20738 29558 20773 29604
rect 20657 29286 20773 29558
rect 20657 29240 20692 29286
rect 20738 29240 20773 29286
rect 20657 28890 20773 29240
rect 21276 29604 21392 29640
rect 21276 29558 21311 29604
rect 21357 29558 21392 29604
rect 21276 29286 21392 29558
rect 21276 29240 21311 29286
rect 21357 29240 21392 29286
rect 21276 28890 21392 29240
rect 21895 29604 22011 29640
rect 21895 29558 21930 29604
rect 21976 29558 22011 29604
rect 21895 29286 22011 29558
rect 21895 29240 21930 29286
rect 21976 29240 22011 29286
rect 21895 28890 22011 29240
rect 22514 29604 22630 29640
rect 22514 29558 22549 29604
rect 22595 29558 22630 29604
rect 22514 29286 22630 29558
rect 22514 29240 22549 29286
rect 22595 29240 22630 29286
rect 22514 28890 22630 29240
rect 230 28725 22630 28890
rect 23082 28962 23760 28986
rect 23082 28924 23369 28962
rect 23421 28924 23760 28962
rect 23082 28878 23211 28924
rect 23257 28878 23369 28924
rect 23421 28910 23527 28924
rect 23415 28878 23527 28910
rect 23573 28878 23760 28924
rect 23082 28776 23760 28878
rect 23082 28724 23369 28776
rect 23421 28724 23760 28776
rect 23082 28703 23760 28724
rect 23082 28587 23230 28703
rect 23082 28541 23143 28587
rect 23189 28541 23230 28587
rect 23082 28405 23230 28541
rect 23082 28359 23143 28405
rect 23189 28359 23230 28405
rect 23082 28224 23230 28359
rect 23082 28178 23143 28224
rect 23189 28178 23230 28224
rect 23082 28042 23230 28178
rect 23082 27996 23143 28042
rect 23189 27996 23230 28042
rect 23082 27811 23230 27996
rect 23335 28587 23450 28623
rect 23335 28541 23369 28587
rect 23415 28541 23450 28587
rect 23335 28405 23450 28541
rect 23335 28359 23369 28405
rect 23415 28372 23450 28405
rect 23335 28224 23386 28359
rect 23335 28178 23369 28224
rect 23438 28216 23450 28372
rect 23415 28178 23450 28216
rect 23335 28042 23450 28178
rect 23335 27996 23369 28042
rect 23415 27996 23450 28042
rect 23335 27959 23450 27996
rect 23555 28587 23760 28703
rect 23555 28541 23679 28587
rect 23725 28541 23760 28587
rect 23555 28405 23760 28541
rect 23555 28359 23679 28405
rect 23725 28359 23760 28405
rect 23555 28224 23760 28359
rect 23555 28178 23679 28224
rect 23725 28178 23760 28224
rect 23555 28042 23760 28178
rect 23555 27996 23679 28042
rect 23725 27996 23760 28042
rect 23082 27765 23143 27811
rect 23189 27765 23230 27811
rect 23082 27630 23230 27765
rect 23082 27584 23143 27630
rect 23189 27584 23230 27630
rect 23082 27449 23230 27584
rect 23082 27403 23143 27449
rect 23189 27403 23230 27449
rect 23082 27267 23230 27403
rect 23082 27221 23143 27267
rect 23189 27221 23230 27267
rect 23082 27184 23230 27221
rect 23335 27811 23450 27848
rect 23335 27765 23369 27811
rect 23415 27765 23450 27811
rect 23335 27630 23450 27765
rect 23335 27593 23369 27630
rect 23335 27437 23347 27593
rect 23415 27584 23450 27630
rect 23399 27449 23450 27584
rect 23335 27403 23369 27437
rect 23415 27403 23450 27449
rect 23335 27267 23450 27403
rect 23335 27221 23369 27267
rect 23415 27221 23450 27267
rect 23335 27184 23450 27221
rect 23555 27811 23760 27996
rect 23555 27765 23679 27811
rect 23725 27765 23760 27811
rect 23555 27630 23760 27765
rect 23555 27584 23679 27630
rect 23725 27584 23760 27630
rect 23555 27449 23760 27584
rect 23555 27403 23679 27449
rect 23725 27403 23760 27449
rect 23555 27267 23760 27403
rect 23555 27221 23679 27267
rect 23725 27221 23760 27267
rect 23555 27184 23760 27221
rect 22263 27031 22913 27105
rect 23249 27093 23624 27104
rect 23249 27047 23328 27093
rect 23468 27047 23624 27093
rect 23249 27030 23624 27047
rect 23259 26943 23305 26956
rect 23259 26835 23305 26897
rect 23259 26727 23305 26789
rect 23259 26619 23305 26681
rect 23259 26511 23305 26573
rect 23259 26417 23305 26465
rect 23144 26405 23305 26417
rect 23144 26249 23156 26405
rect 23208 26403 23305 26405
rect 23208 26357 23259 26403
rect 23208 26295 23305 26357
rect 23208 26249 23259 26295
rect 23144 26237 23305 26249
rect 23259 26188 23305 26237
rect 23259 26081 23305 26142
rect 23259 25974 23305 26035
rect 23259 25867 23305 25928
rect 23259 25760 23305 25821
rect 23259 25653 23305 25714
rect 23259 25594 23305 25607
rect 23483 26943 23529 26956
rect 23483 26835 23529 26897
rect 23483 26727 23529 26789
rect 23483 26619 23529 26681
rect 23483 26511 23529 26573
rect 23483 26417 23529 26465
rect 23483 26405 23644 26417
rect 23483 26403 23580 26405
rect 23529 26357 23580 26403
rect 23483 26295 23580 26357
rect 23529 26249 23580 26295
rect 23632 26249 23644 26405
rect 23483 26237 23644 26249
rect 23483 26188 23529 26237
rect 23483 26081 23529 26142
rect 23483 25974 23529 26035
rect 23483 25867 23529 25928
rect 23483 25760 23529 25821
rect 23483 25653 23529 25714
rect 23483 25594 23529 25607
rect 23153 25357 23635 25369
rect 23153 25356 23571 25357
rect 23153 25310 23257 25356
rect 23303 25310 23481 25356
rect 23527 25310 23571 25356
rect 23153 25248 23571 25310
rect 23153 25202 23257 25248
rect 23303 25202 23481 25248
rect 23527 25202 23571 25248
rect 23153 25201 23571 25202
rect 23623 25201 23635 25357
rect 23153 25189 23635 25201
rect 23153 25140 23632 25189
rect 23153 25094 23257 25140
rect 23303 25094 23481 25140
rect 23527 25094 23632 25140
rect 23153 25032 23632 25094
rect 23153 24986 23257 25032
rect 23303 24986 23481 25032
rect 23527 24986 23632 25032
rect 23153 24924 23632 24986
rect 23153 24878 23257 24924
rect 23303 24878 23481 24924
rect 23527 24878 23632 24924
rect 23153 24816 23632 24878
rect 23153 24770 23257 24816
rect 23303 24770 23481 24816
rect 23527 24770 23632 24816
rect 23153 24708 23632 24770
rect 23153 24662 23257 24708
rect 23303 24662 23481 24708
rect 23527 24662 23632 24708
rect 23153 24601 23632 24662
rect 23153 24555 23257 24601
rect 23303 24555 23481 24601
rect 23527 24555 23632 24601
rect 23153 24494 23632 24555
rect 23153 24448 23257 24494
rect 23303 24448 23481 24494
rect 23527 24448 23632 24494
rect 23153 24387 23632 24448
rect 23153 24341 23257 24387
rect 23303 24341 23481 24387
rect 23527 24341 23632 24387
rect 23153 24280 23632 24341
rect 23153 24234 23257 24280
rect 23303 24234 23481 24280
rect 23527 24234 23632 24280
rect 23153 24173 23632 24234
rect 23153 24127 23257 24173
rect 23303 24127 23481 24173
rect 23527 24127 23632 24173
rect 23153 24066 23632 24127
rect 23153 24020 23257 24066
rect 23303 24020 23481 24066
rect 23527 24020 23632 24066
rect 23153 24007 23632 24020
rect 23153 23678 23223 24007
rect 23302 23926 23483 23937
rect 23302 23922 23369 23926
rect 23302 23766 23349 23922
rect 23415 23880 23483 23926
rect 23401 23766 23483 23880
rect 23302 23754 23483 23766
rect 23561 23678 23632 24007
rect 23153 23665 23303 23678
rect 23153 23619 23257 23665
rect 23153 23557 23303 23619
rect 23153 23511 23257 23557
rect 23153 23449 23303 23511
rect 23153 23403 23257 23449
rect 23153 23341 23303 23403
rect 23153 23295 23257 23341
rect 23153 23233 23303 23295
rect 23153 23187 23257 23233
rect 23153 23125 23303 23187
rect 23153 23079 23257 23125
rect 23153 23017 23303 23079
rect 23153 22971 23257 23017
rect 23153 22910 23303 22971
rect 23153 22864 23257 22910
rect 23153 22803 23303 22864
rect 23153 22757 23257 22803
rect 23153 22696 23303 22757
rect 23153 22650 23257 22696
rect 23153 22589 23303 22650
rect 23153 22543 23257 22589
rect 23153 22482 23303 22543
rect 23153 22436 23257 22482
rect 23153 22416 23303 22436
rect 23481 23665 23632 23678
rect 23527 23619 23632 23665
rect 23481 23557 23632 23619
rect 23527 23511 23632 23557
rect 23481 23449 23632 23511
rect 23527 23403 23632 23449
rect 23481 23341 23632 23403
rect 23527 23295 23632 23341
rect 23481 23233 23632 23295
rect 23527 23187 23632 23233
rect 23481 23125 23632 23187
rect 23527 23079 23632 23125
rect 23481 23017 23632 23079
rect 23527 22971 23632 23017
rect 23481 22910 23632 22971
rect 23527 22864 23632 22910
rect 23481 22803 23632 22864
rect 23527 22757 23632 22803
rect 23481 22696 23632 22757
rect 23527 22650 23632 22696
rect 23481 22589 23632 22650
rect 23527 22543 23632 22589
rect 23481 22482 23632 22543
rect 23527 22436 23632 22482
rect 23153 22375 23338 22416
rect 23153 22329 23257 22375
rect 23303 22329 23338 22375
rect 23153 22326 23338 22329
rect 23245 22246 23338 22326
rect 23481 22375 23632 22436
rect 23527 22329 23632 22375
rect 23481 22316 23632 22329
rect 23245 22242 23657 22246
rect 23245 22222 23856 22242
rect 23245 22170 23578 22222
rect 23630 22170 23764 22222
rect 23816 22170 23856 22222
rect 23245 22150 23856 22170
rect 23245 22149 23657 22150
rect 23631 22065 23773 22070
rect 23082 22024 23773 22065
rect 23082 21972 23536 22024
rect 23588 22019 23773 22024
rect 23588 21973 23679 22019
rect 23725 21973 23773 22019
rect 23588 21972 23773 21973
rect 23082 21931 23773 21972
rect 23631 21922 23773 21931
rect 23141 21820 23654 21843
rect 23141 21768 23156 21820
rect 23208 21768 23654 21820
rect 23141 21746 23654 21768
rect 23561 21674 23654 21746
rect 23153 21661 23303 21674
rect 23153 21615 23257 21661
rect 23153 21553 23303 21615
rect 23153 21507 23257 21553
rect 23153 21445 23303 21507
rect 23153 21399 23257 21445
rect 23153 21337 23303 21399
rect 23153 21291 23257 21337
rect 23153 21229 23303 21291
rect 23153 21183 23257 21229
rect 23153 21121 23303 21183
rect 23153 21075 23257 21121
rect 23153 21013 23303 21075
rect 23153 20967 23257 21013
rect 23153 20906 23303 20967
rect 23153 20860 23257 20906
rect 23153 20799 23303 20860
rect 23153 20753 23257 20799
rect 23153 20692 23303 20753
rect 23153 20646 23257 20692
rect 23153 20585 23303 20646
rect 23153 20539 23257 20585
rect 23153 20478 23303 20539
rect 23153 20432 23257 20478
rect 23153 20371 23303 20432
rect 23153 20325 23257 20371
rect 23153 20312 23303 20325
rect 23481 21661 23654 21674
rect 23527 21615 23654 21661
rect 23481 21553 23654 21615
rect 23527 21507 23654 21553
rect 23481 21445 23654 21507
rect 23527 21399 23654 21445
rect 23481 21337 23654 21399
rect 23527 21291 23654 21337
rect 23481 21229 23654 21291
rect 23527 21183 23654 21229
rect 23481 21121 23654 21183
rect 23527 21075 23654 21121
rect 23481 21013 23654 21075
rect 23527 20967 23654 21013
rect 23481 20906 23654 20967
rect 23527 20860 23654 20906
rect 23481 20799 23654 20860
rect 23527 20753 23654 20799
rect 23481 20692 23654 20753
rect 23527 20646 23654 20692
rect 23481 20585 23654 20646
rect 23527 20539 23654 20585
rect 23481 20478 23654 20539
rect 23527 20432 23654 20478
rect 23481 20371 23654 20432
rect 23527 20325 23654 20371
rect 23481 20312 23654 20325
rect 23153 19819 23223 20312
rect 23302 20228 23483 20242
rect 23302 20182 23369 20228
rect 23415 20182 23483 20228
rect 23302 20179 23483 20182
rect 23302 20127 23364 20179
rect 23416 20127 23483 20179
rect 23302 20107 23483 20127
rect 23302 19984 23483 20027
rect 23302 19932 23314 19984
rect 23470 19932 23483 19984
rect 23302 19905 23369 19932
rect 23415 19905 23483 19932
rect 23302 19891 23483 19905
rect 23561 19819 23654 20312
rect 23153 19818 23303 19819
rect 23481 19818 23654 19819
rect 23153 19806 23654 19818
rect 23153 19760 23257 19806
rect 23303 19760 23481 19806
rect 23527 19760 23654 19806
rect 23153 19698 23654 19760
rect 23153 19652 23257 19698
rect 23303 19652 23481 19698
rect 23527 19652 23654 19698
rect 23153 19590 23654 19652
rect 23153 19544 23257 19590
rect 23303 19544 23481 19590
rect 23527 19544 23654 19590
rect 23153 19482 23654 19544
rect 23153 19436 23257 19482
rect 23303 19436 23481 19482
rect 23527 19436 23654 19482
rect 23153 19374 23654 19436
rect 23153 19328 23257 19374
rect 23303 19328 23481 19374
rect 23527 19328 23654 19374
rect 23153 19266 23654 19328
rect 23153 19220 23257 19266
rect 23303 19220 23481 19266
rect 23527 19220 23654 19266
rect 23153 19158 23654 19220
rect 23153 19112 23257 19158
rect 23303 19112 23481 19158
rect 23527 19112 23654 19158
rect 23153 19051 23654 19112
rect 23153 19005 23257 19051
rect 23303 19005 23481 19051
rect 23527 19005 23654 19051
rect 23153 18944 23654 19005
rect 23153 18898 23257 18944
rect 23303 18898 23481 18944
rect 23527 18898 23654 18944
rect 23153 18837 23654 18898
rect 23153 18791 23257 18837
rect 23303 18791 23481 18837
rect 23527 18791 23654 18837
rect 23153 18730 23654 18791
rect 23153 18684 23257 18730
rect 23303 18684 23481 18730
rect 23527 18684 23654 18730
rect 23153 18623 23654 18684
rect 23153 18577 23257 18623
rect 23303 18577 23481 18623
rect 23527 18577 23654 18623
rect 23153 18516 23654 18577
rect 23153 18470 23257 18516
rect 23303 18470 23481 18516
rect 23527 18470 23654 18516
rect 23153 18467 23654 18470
rect 23153 18457 23552 18467
rect 23153 18433 23338 18457
rect 22779 18313 23338 18433
rect 22779 16586 22895 18313
rect 23082 18183 23760 18211
rect 23082 18131 23139 18183
rect 23191 18174 23319 18183
rect 23371 18174 23760 18183
rect 23191 18131 23205 18174
rect 23082 18128 23205 18131
rect 23251 18131 23319 18174
rect 23251 18128 23363 18131
rect 23409 18128 23521 18174
rect 23567 18128 23679 18174
rect 23725 18128 23760 18174
rect 23082 18091 23760 18128
rect 23082 17835 23153 18091
rect 23518 18011 23760 18091
rect 23257 17988 23760 18011
rect 23257 17936 23295 17988
rect 23347 17984 23760 17988
rect 23347 17938 23426 17984
rect 23472 17938 23760 17984
rect 23347 17936 23760 17938
rect 23257 17914 23760 17936
rect 23082 17719 23256 17835
rect 23082 17673 23176 17719
rect 23222 17673 23256 17719
rect 23082 17556 23256 17673
rect 23379 17823 23507 17835
rect 23379 17719 23443 17823
rect 23379 17673 23426 17719
rect 23379 17667 23443 17673
rect 23495 17667 23507 17823
rect 23379 17556 23507 17667
rect 23645 17719 23759 17914
rect 23645 17673 23679 17719
rect 23725 17673 23759 17719
rect 23645 17556 23759 17673
rect 23082 17222 23263 17259
rect 23082 17176 23217 17222
rect 23082 17030 23263 17176
rect 23414 17222 23487 17556
rect 23414 17176 23441 17222
rect 23414 17139 23487 17176
rect 23645 17222 23760 17259
rect 23645 17176 23665 17222
rect 23711 17176 23760 17222
rect 23645 17030 23760 17176
rect 23082 16939 23760 17030
rect 23082 16923 23366 16939
rect 23418 16923 23760 16939
rect 23082 16877 23247 16923
rect 23669 16877 23760 16923
rect 23082 16835 23760 16877
rect 22779 16466 23910 16586
rect 23141 15609 23573 15645
rect 23141 15608 23216 15609
rect 23268 15608 23402 15609
rect 23141 15562 23176 15608
rect 23268 15562 23334 15608
rect 23380 15562 23402 15608
rect 23141 15557 23216 15562
rect 23268 15557 23402 15562
rect 23454 15608 23573 15609
rect 23454 15562 23492 15608
rect 23538 15562 23573 15608
rect 23454 15557 23573 15562
rect 23141 15525 23573 15557
rect 23168 15158 23214 15171
rect 23168 15053 23214 15112
rect 23144 15015 23168 15045
rect 23392 15158 23438 15171
rect 23392 15053 23438 15112
rect 23214 15015 23236 15045
rect 23144 14963 23164 15015
rect 23216 14963 23236 15015
rect 23144 14948 23236 14963
rect 23144 14902 23168 14948
rect 23214 14902 23236 14948
rect 23144 14843 23236 14902
rect 23144 14829 23168 14843
rect 23214 14829 23236 14843
rect 23144 14777 23164 14829
rect 23216 14777 23236 14829
rect 23616 15158 23662 15171
rect 23616 15053 23662 15112
rect 23392 14948 23438 15007
rect 23392 14843 23438 14902
rect 23392 14783 23438 14797
rect 23592 15015 23616 15045
rect 23662 15015 23684 15045
rect 23592 14963 23612 15015
rect 23664 14963 23684 15015
rect 23592 14948 23684 14963
rect 23592 14902 23616 14948
rect 23662 14902 23684 14948
rect 23592 14843 23684 14902
rect 23592 14829 23616 14843
rect 23662 14829 23684 14843
rect 23144 14738 23236 14777
rect 23144 14737 23168 14738
rect 23214 14737 23236 14738
rect 23356 14738 23473 14783
rect 23168 14633 23214 14692
rect 23168 14528 23214 14587
rect 23168 14469 23214 14482
rect 23356 14692 23392 14738
rect 23438 14692 23473 14738
rect 23592 14777 23612 14829
rect 23664 14777 23684 14829
rect 23592 14738 23684 14777
rect 23592 14737 23616 14738
rect 23356 14633 23473 14692
rect 23356 14587 23392 14633
rect 23438 14587 23473 14633
rect 23356 14528 23473 14587
rect 23356 14482 23392 14528
rect 23438 14482 23473 14528
rect 23356 14398 23473 14482
rect 23662 14737 23684 14738
rect 23616 14633 23662 14692
rect 23616 14528 23662 14587
rect 23616 14469 23662 14482
rect 22955 14323 23473 14398
rect 23793 14384 23910 16466
rect 22955 10723 23027 14323
rect 23168 14152 23214 14165
rect 23132 13902 23168 13938
rect 23356 14152 23473 14323
rect 23563 14347 23910 14384
rect 23563 14301 23598 14347
rect 23644 14301 23756 14347
rect 23802 14301 23910 14347
rect 23563 14264 23910 14301
rect 23356 14060 23392 14152
rect 23214 13902 23249 13938
rect 23132 13664 23249 13902
rect 23438 14060 23473 14152
rect 23616 14152 23662 14165
rect 23392 13889 23438 13902
rect 23580 13902 23616 13938
rect 23662 13902 23697 13938
rect 23580 13664 23697 13902
rect 23132 13613 23697 13664
rect 23132 13567 23233 13613
rect 23279 13567 23391 13613
rect 23437 13567 23549 13613
rect 23595 13567 23697 13613
rect 23132 13516 23697 13567
rect 23132 12576 23249 13516
rect 23132 12524 23169 12576
rect 23221 12524 23249 12576
rect 23132 12491 23249 12524
rect 23132 12390 23172 12491
rect 23218 12390 23249 12491
rect 23132 12338 23169 12390
rect 23221 12338 23249 12390
rect 23132 12038 23172 12338
rect 23218 12038 23249 12338
rect 23132 11986 23169 12038
rect 23221 11986 23249 12038
rect 23132 11852 23172 11986
rect 23218 11852 23249 11986
rect 23132 11800 23169 11852
rect 23221 11800 23249 11852
rect 23132 11719 23172 11800
rect 23149 11433 23172 11463
rect 23218 11719 23249 11800
rect 23356 12576 23486 12616
rect 23356 12524 23395 12576
rect 23447 12524 23486 12576
rect 23356 12491 23486 12524
rect 23356 12358 23396 12491
rect 23442 12358 23486 12491
rect 23356 12306 23395 12358
rect 23447 12306 23486 12358
rect 23356 12140 23396 12306
rect 23442 12140 23486 12306
rect 23356 12088 23395 12140
rect 23447 12088 23486 12140
rect 23356 11923 23396 12088
rect 23442 11923 23486 12088
rect 23356 11871 23395 11923
rect 23447 11871 23486 11923
rect 23356 11705 23396 11871
rect 23442 11705 23486 11871
rect 23580 12576 23697 13516
rect 23580 12524 23610 12576
rect 23662 12524 23697 12576
rect 23580 12491 23697 12524
rect 23580 12390 23620 12491
rect 23580 12338 23610 12390
rect 23580 12038 23620 12338
rect 23580 11986 23610 12038
rect 23580 11852 23620 11986
rect 23580 11800 23610 11852
rect 23580 11719 23620 11800
rect 23356 11653 23395 11705
rect 23447 11653 23486 11705
rect 23356 11487 23396 11653
rect 23442 11487 23486 11653
rect 23218 11433 23241 11463
rect 23149 11381 23169 11433
rect 23221 11381 23241 11433
rect 23149 11247 23172 11381
rect 23218 11247 23241 11381
rect 23149 11195 23169 11247
rect 23221 11195 23241 11247
rect 23149 11155 23172 11195
rect 23218 11155 23241 11195
rect 23356 11435 23395 11487
rect 23447 11435 23486 11487
rect 23356 11270 23396 11435
rect 23442 11270 23486 11435
rect 23356 11218 23395 11270
rect 23447 11218 23486 11270
rect 23172 10804 23218 10817
rect 23356 11052 23396 11218
rect 23442 11052 23486 11218
rect 23590 11433 23620 11463
rect 23666 11719 23697 12491
rect 23590 11381 23610 11433
rect 23590 11247 23620 11381
rect 23590 11195 23610 11247
rect 23590 11155 23620 11195
rect 23356 11000 23395 11052
rect 23447 11000 23486 11052
rect 23356 10835 23396 11000
rect 23442 10835 23486 11000
rect 23356 10783 23395 10835
rect 23447 10783 23486 10835
rect 23666 11155 23682 11463
rect 23620 10804 23666 10817
rect 22955 10686 23253 10723
rect 22955 10640 23014 10686
rect 23060 10640 23172 10686
rect 23218 10640 23253 10686
rect 22955 10603 23253 10640
rect 23356 10617 23486 10783
rect 23356 10565 23395 10617
rect 23447 10565 23486 10617
rect 23172 10510 23218 10523
rect 23172 10407 23218 10464
rect 23172 10304 23218 10361
rect 23172 10201 23218 10258
rect 23172 10098 23218 10155
rect 23172 9995 23218 10052
rect 23172 9892 23218 9949
rect 23172 9789 23218 9846
rect 23172 9686 23218 9743
rect 23172 9583 23218 9640
rect 23172 9480 23218 9537
rect 23172 9377 23218 9434
rect 23172 9274 23218 9331
rect 23172 9171 23218 9228
rect 23172 9068 23218 9125
rect 23172 8965 23218 9022
rect 23172 8862 23218 8919
rect 23137 8408 23172 8519
rect 23356 10510 23486 10565
rect 23356 10464 23396 10510
rect 23442 10464 23486 10510
rect 23356 10407 23486 10464
rect 23356 10399 23396 10407
rect 23442 10399 23486 10407
rect 23356 10347 23395 10399
rect 23447 10347 23486 10399
rect 23356 10304 23486 10347
rect 23356 10258 23396 10304
rect 23442 10258 23486 10304
rect 23356 10201 23486 10258
rect 23356 10182 23396 10201
rect 23442 10182 23486 10201
rect 23356 10130 23395 10182
rect 23447 10130 23486 10182
rect 23356 10098 23486 10130
rect 23356 10052 23396 10098
rect 23442 10052 23486 10098
rect 23356 9995 23486 10052
rect 23356 9964 23396 9995
rect 23442 9964 23486 9995
rect 23356 9912 23395 9964
rect 23447 9912 23486 9964
rect 23356 9892 23486 9912
rect 23356 9846 23396 9892
rect 23442 9846 23486 9892
rect 23356 9789 23486 9846
rect 23356 9746 23396 9789
rect 23442 9746 23486 9789
rect 23356 9694 23395 9746
rect 23447 9694 23486 9746
rect 23356 9686 23486 9694
rect 23356 9640 23396 9686
rect 23442 9640 23486 9686
rect 23356 9583 23486 9640
rect 23356 9537 23396 9583
rect 23442 9537 23486 9583
rect 23356 9529 23486 9537
rect 23356 9477 23395 9529
rect 23447 9477 23486 9529
rect 23356 9434 23396 9477
rect 23442 9434 23486 9477
rect 23356 9377 23486 9434
rect 23356 9331 23396 9377
rect 23442 9331 23486 9377
rect 23356 9311 23486 9331
rect 23356 9259 23395 9311
rect 23447 9259 23486 9311
rect 23356 9228 23396 9259
rect 23442 9228 23486 9259
rect 23356 9171 23486 9228
rect 23356 9125 23396 9171
rect 23442 9125 23486 9171
rect 23356 9093 23486 9125
rect 23356 9041 23395 9093
rect 23447 9041 23486 9093
rect 23356 9022 23396 9041
rect 23442 9022 23486 9041
rect 23356 8965 23486 9022
rect 23356 8919 23396 8965
rect 23442 8919 23486 8965
rect 23356 8876 23486 8919
rect 23356 8824 23395 8876
rect 23447 8824 23486 8876
rect 23356 8658 23396 8824
rect 23442 8658 23486 8824
rect 23356 8606 23395 8658
rect 23447 8606 23486 8658
rect 23218 8408 23253 8519
rect 23137 7774 23253 8408
rect 23137 7722 23173 7774
rect 23225 7722 23253 7774
rect 23137 7588 23253 7722
rect 23137 7536 23173 7588
rect 23225 7536 23253 7588
rect 23137 7402 23253 7536
rect 23137 7350 23173 7402
rect 23225 7350 23253 7402
rect 23137 7325 23253 7350
rect 23024 7288 23253 7325
rect 23024 7242 23058 7288
rect 23104 7242 23253 7288
rect 23024 7205 23253 7242
rect 23356 8441 23396 8606
rect 23442 8441 23486 8606
rect 23620 10510 23666 10523
rect 23620 10407 23666 10464
rect 23620 10304 23666 10361
rect 23620 10201 23666 10258
rect 23620 10098 23666 10155
rect 23620 9995 23666 10052
rect 23620 9892 23666 9949
rect 23620 9789 23666 9846
rect 23620 9686 23666 9743
rect 23620 9583 23666 9640
rect 23620 9480 23666 9537
rect 23620 9377 23666 9434
rect 23620 9274 23666 9331
rect 23620 9171 23666 9228
rect 23620 9068 23666 9125
rect 23620 8965 23666 9022
rect 23620 8862 23666 8919
rect 23356 8389 23395 8441
rect 23447 8389 23486 8441
rect 23356 8223 23486 8389
rect 23356 8171 23395 8223
rect 23447 8171 23486 8223
rect 23356 8005 23486 8171
rect 23356 7953 23395 8005
rect 23447 7953 23486 8005
rect 23356 7788 23486 7953
rect 23356 7736 23395 7788
rect 23447 7736 23486 7788
rect 23356 7570 23486 7736
rect 23356 7518 23395 7570
rect 23447 7518 23486 7570
rect 23356 7352 23486 7518
rect 23356 7300 23395 7352
rect 23447 7300 23486 7352
rect 23585 8408 23620 8519
rect 23666 8408 23701 8519
rect 23585 7774 23701 8408
rect 23585 7722 23615 7774
rect 23667 7722 23701 7774
rect 23585 7588 23701 7722
rect 23585 7536 23615 7588
rect 23667 7536 23701 7588
rect 23585 7402 23701 7536
rect 23585 7350 23615 7402
rect 23667 7350 23701 7402
rect 23585 7325 23701 7350
rect 23356 7042 23486 7300
rect 23568 7288 23701 7325
rect 23568 7242 23602 7288
rect 23648 7242 23701 7288
rect 23568 7205 23701 7242
rect 23308 5013 23530 7042
rect 23259 4973 23599 5013
rect 23259 4921 23297 4973
rect 23349 4921 23509 4973
rect 23561 4921 23599 4973
rect 23259 4755 23599 4921
rect 23259 4703 23297 4755
rect 23349 4703 23509 4755
rect 23561 4703 23599 4755
rect 23259 4662 23599 4703
<< via1 >>
rect 66 89396 69 89535
rect 69 89396 115 89535
rect 115 89396 118 89535
rect 66 89275 118 89396
rect 23894 89472 23946 89477
rect 23894 89426 23899 89472
rect 23899 89426 23945 89472
rect 23945 89426 23946 89472
rect 23894 89425 23946 89426
rect 23894 89207 23946 89259
rect 66 87877 118 87936
rect 66 87737 69 87877
rect 69 87737 115 87877
rect 115 87737 118 87877
rect 66 87676 118 87737
rect 23894 87912 23946 87940
rect 23894 87888 23899 87912
rect 23899 87888 23945 87912
rect 23945 87888 23946 87912
rect 23894 87702 23899 87722
rect 23899 87702 23945 87722
rect 23945 87702 23946 87722
rect 23894 87670 23946 87702
rect 66 86077 118 86137
rect 66 85937 69 86077
rect 69 85937 115 86077
rect 115 85937 118 86077
rect 66 85877 118 85937
rect 23894 86112 23946 86140
rect 23894 86088 23899 86112
rect 23899 86088 23945 86112
rect 23945 86088 23946 86112
rect 23894 85902 23899 85922
rect 23899 85902 23945 85922
rect 23945 85902 23946 85922
rect 23894 85870 23946 85902
rect 66 84277 118 84337
rect 66 84137 69 84277
rect 69 84137 115 84277
rect 115 84137 118 84277
rect 66 84077 118 84137
rect 23894 84312 23946 84340
rect 23894 84288 23899 84312
rect 23899 84288 23945 84312
rect 23945 84288 23946 84312
rect 23894 84102 23899 84122
rect 23899 84102 23945 84122
rect 23945 84102 23946 84122
rect 23894 84070 23946 84102
rect 66 82477 118 82537
rect 66 82337 69 82477
rect 69 82337 115 82477
rect 115 82337 118 82477
rect 66 82277 118 82337
rect 23894 82512 23946 82540
rect 23894 82488 23899 82512
rect 23899 82488 23945 82512
rect 23945 82488 23946 82512
rect 23894 82302 23899 82322
rect 23899 82302 23945 82322
rect 23945 82302 23946 82322
rect 23894 82270 23946 82302
rect 66 80677 118 80736
rect 66 80537 69 80677
rect 69 80537 115 80677
rect 115 80537 118 80677
rect 66 80476 118 80537
rect 23894 80712 23946 80740
rect 23894 80688 23899 80712
rect 23899 80688 23945 80712
rect 23945 80688 23946 80712
rect 23894 80502 23899 80522
rect 23899 80502 23945 80522
rect 23945 80502 23946 80522
rect 23894 80470 23946 80502
rect 66 78877 118 78937
rect 66 78737 69 78877
rect 69 78737 115 78877
rect 115 78737 118 78877
rect 66 78677 118 78737
rect 23894 78912 23946 78940
rect 23894 78888 23899 78912
rect 23899 78888 23945 78912
rect 23945 78888 23946 78912
rect 23894 78702 23899 78722
rect 23899 78702 23945 78722
rect 23945 78702 23946 78722
rect 23894 78670 23946 78702
rect 66 77077 118 77138
rect 66 76937 69 77077
rect 69 76937 115 77077
rect 115 76937 118 77077
rect 66 76878 118 76937
rect 23894 77112 23946 77140
rect 23894 77088 23899 77112
rect 23899 77088 23945 77112
rect 23945 77088 23946 77112
rect 23894 76902 23899 76922
rect 23899 76902 23945 76922
rect 23945 76902 23946 76922
rect 23894 76870 23946 76902
rect 66 75277 118 75337
rect 66 75137 69 75277
rect 69 75137 115 75277
rect 115 75137 118 75277
rect 66 75077 118 75137
rect 23894 75312 23946 75340
rect 23894 75288 23899 75312
rect 23899 75288 23945 75312
rect 23945 75288 23946 75312
rect 23894 75102 23899 75122
rect 23899 75102 23945 75122
rect 23945 75102 23946 75122
rect 23894 75070 23946 75102
rect 66 73477 118 73537
rect 66 73337 69 73477
rect 69 73337 115 73477
rect 115 73337 118 73477
rect 66 73277 118 73337
rect 23894 73512 23946 73540
rect 23894 73488 23899 73512
rect 23899 73488 23945 73512
rect 23945 73488 23946 73512
rect 23894 73302 23899 73322
rect 23899 73302 23945 73322
rect 23945 73302 23946 73322
rect 23894 73270 23946 73302
rect 66 71677 118 71737
rect 66 71537 69 71677
rect 69 71537 115 71677
rect 115 71537 118 71677
rect 66 71477 118 71537
rect 23894 71712 23946 71740
rect 23894 71688 23899 71712
rect 23899 71688 23945 71712
rect 23945 71688 23946 71712
rect 23894 71502 23899 71522
rect 23899 71502 23945 71522
rect 23945 71502 23946 71522
rect 23894 71470 23946 71502
rect 66 69877 118 69937
rect 66 69737 69 69877
rect 69 69737 115 69877
rect 115 69737 118 69877
rect 66 69677 118 69737
rect 23894 69912 23946 69940
rect 23894 69888 23899 69912
rect 23899 69888 23945 69912
rect 23945 69888 23946 69912
rect 23894 69702 23899 69722
rect 23899 69702 23945 69722
rect 23945 69702 23946 69722
rect 23894 69670 23946 69702
rect 66 68077 118 68137
rect 66 67937 69 68077
rect 69 67937 115 68077
rect 115 67937 118 68077
rect 66 67877 118 67937
rect 23894 68112 23946 68140
rect 23894 68088 23899 68112
rect 23899 68088 23945 68112
rect 23945 68088 23946 68112
rect 23894 67902 23899 67922
rect 23899 67902 23945 67922
rect 23945 67902 23946 67922
rect 23894 67870 23946 67902
rect 66 66277 118 66337
rect 66 66137 69 66277
rect 69 66137 115 66277
rect 115 66137 118 66277
rect 66 66077 118 66137
rect 23894 66312 23946 66340
rect 23894 66288 23899 66312
rect 23899 66288 23945 66312
rect 23945 66288 23946 66312
rect 23894 66102 23899 66122
rect 23899 66102 23945 66122
rect 23945 66102 23946 66122
rect 23894 66070 23946 66102
rect 66 64477 118 64537
rect 66 64337 69 64477
rect 69 64337 115 64477
rect 115 64337 118 64477
rect 66 64277 118 64337
rect 23894 64512 23946 64540
rect 23894 64488 23899 64512
rect 23899 64488 23945 64512
rect 23945 64488 23946 64512
rect 23894 64302 23899 64322
rect 23899 64302 23945 64322
rect 23945 64302 23946 64322
rect 23894 64270 23946 64302
rect 66 62677 118 62737
rect 66 62537 69 62677
rect 69 62537 115 62677
rect 115 62537 118 62677
rect 66 62477 118 62537
rect 23894 62712 23946 62740
rect 23894 62688 23899 62712
rect 23899 62688 23945 62712
rect 23945 62688 23946 62712
rect 23894 62502 23899 62522
rect 23899 62502 23945 62522
rect 23945 62502 23946 62522
rect 23894 62470 23946 62502
rect 66 60877 118 60937
rect 66 60737 69 60877
rect 69 60737 115 60877
rect 115 60737 118 60877
rect 66 60677 118 60737
rect 23894 60912 23946 60940
rect 23894 60888 23899 60912
rect 23899 60888 23945 60912
rect 23945 60888 23946 60912
rect 23894 60702 23899 60722
rect 23899 60702 23945 60722
rect 23945 60702 23946 60722
rect 23894 60670 23946 60702
rect 66 59077 118 59137
rect 66 58937 69 59077
rect 69 58937 115 59077
rect 115 58937 118 59077
rect 66 58877 118 58937
rect 23894 59112 23946 59140
rect 23894 59088 23899 59112
rect 23899 59088 23945 59112
rect 23945 59088 23946 59112
rect 23894 58902 23899 58922
rect 23899 58902 23945 58922
rect 23945 58902 23946 58922
rect 23894 58870 23946 58902
rect 66 57277 118 57337
rect 66 57137 69 57277
rect 69 57137 115 57277
rect 115 57137 118 57277
rect 66 57077 118 57137
rect 23894 57312 23946 57340
rect 23894 57288 23899 57312
rect 23899 57288 23945 57312
rect 23945 57288 23946 57312
rect 23894 57102 23899 57122
rect 23899 57102 23945 57122
rect 23945 57102 23946 57122
rect 23894 57070 23946 57102
rect 66 55477 118 55537
rect 66 55337 69 55477
rect 69 55337 115 55477
rect 115 55337 118 55477
rect 66 55277 118 55337
rect 23894 55512 23946 55544
rect 23894 55492 23899 55512
rect 23899 55492 23945 55512
rect 23945 55492 23946 55512
rect 23894 55302 23899 55326
rect 23899 55302 23945 55326
rect 23945 55302 23946 55326
rect 23894 55274 23946 55302
rect 62 53677 114 53737
rect 62 53537 69 53677
rect 69 53537 114 53677
rect 62 53477 114 53537
rect 23894 53712 23946 53740
rect 23894 53688 23899 53712
rect 23899 53688 23945 53712
rect 23945 53688 23946 53712
rect 23894 53502 23899 53522
rect 23899 53502 23945 53522
rect 23945 53502 23946 53522
rect 23894 53470 23946 53502
rect 66 51877 118 51937
rect 66 51737 69 51877
rect 69 51737 115 51877
rect 115 51737 118 51877
rect 66 51677 118 51737
rect 23894 51912 23946 51944
rect 23894 51892 23899 51912
rect 23899 51892 23945 51912
rect 23945 51892 23946 51912
rect 23894 51702 23899 51726
rect 23899 51702 23945 51726
rect 23945 51702 23946 51726
rect 23894 51674 23946 51702
rect 66 50077 118 50137
rect 66 49937 69 50077
rect 69 49937 115 50077
rect 115 49937 118 50077
rect 66 49877 118 49937
rect 23894 50112 23946 50140
rect 23894 50088 23899 50112
rect 23899 50088 23945 50112
rect 23945 50088 23946 50112
rect 23894 49902 23899 49922
rect 23899 49902 23945 49922
rect 23945 49902 23946 49922
rect 23894 49870 23946 49902
rect 66 48277 118 48337
rect 66 48137 69 48277
rect 69 48137 115 48277
rect 115 48137 118 48277
rect 66 48077 118 48137
rect 23894 48312 23946 48344
rect 23894 48292 23899 48312
rect 23899 48292 23945 48312
rect 23945 48292 23946 48312
rect 23894 48102 23899 48126
rect 23899 48102 23945 48126
rect 23945 48102 23946 48126
rect 23894 48074 23946 48102
rect 66 46477 118 46537
rect 66 46337 69 46477
rect 69 46337 115 46477
rect 115 46337 118 46477
rect 66 46277 118 46337
rect 23894 46512 23946 46540
rect 23894 46488 23899 46512
rect 23899 46488 23945 46512
rect 23945 46488 23946 46512
rect 23894 46302 23899 46322
rect 23899 46302 23945 46322
rect 23945 46302 23946 46322
rect 23894 46270 23946 46302
rect 66 44677 118 44737
rect 66 44537 69 44677
rect 69 44537 115 44677
rect 115 44537 118 44677
rect 66 44477 118 44537
rect 23894 44712 23946 44744
rect 23894 44692 23899 44712
rect 23899 44692 23945 44712
rect 23945 44692 23946 44712
rect 23894 44502 23899 44526
rect 23899 44502 23945 44526
rect 23945 44502 23946 44526
rect 23894 44474 23946 44502
rect 66 42877 118 42937
rect 66 42737 69 42877
rect 69 42737 115 42877
rect 115 42737 118 42877
rect 66 42677 118 42737
rect 23894 42912 23946 42940
rect 23894 42888 23899 42912
rect 23899 42888 23945 42912
rect 23945 42888 23946 42912
rect 23894 42702 23899 42722
rect 23899 42702 23945 42722
rect 23945 42702 23946 42722
rect 23894 42670 23946 42702
rect 66 41077 118 41137
rect 66 40937 69 41077
rect 69 40937 115 41077
rect 115 40937 118 41077
rect 66 40877 118 40937
rect 23894 41112 23946 41144
rect 23894 41092 23899 41112
rect 23899 41092 23945 41112
rect 23945 41092 23946 41112
rect 23894 40902 23899 40926
rect 23899 40902 23945 40926
rect 23945 40902 23946 40926
rect 23894 40874 23946 40902
rect 66 39277 118 39337
rect 66 39137 69 39277
rect 69 39137 115 39277
rect 115 39137 118 39277
rect 66 39077 118 39137
rect 23894 39312 23946 39340
rect 23894 39288 23899 39312
rect 23899 39288 23945 39312
rect 23945 39288 23946 39312
rect 23894 39102 23899 39122
rect 23899 39102 23945 39122
rect 23945 39102 23946 39122
rect 23894 39070 23946 39102
rect 66 37477 118 37537
rect 66 37337 69 37477
rect 69 37337 115 37477
rect 115 37337 118 37477
rect 66 37277 118 37337
rect 23894 37512 23946 37544
rect 23894 37492 23899 37512
rect 23899 37492 23945 37512
rect 23945 37492 23946 37512
rect 23894 37302 23899 37326
rect 23899 37302 23945 37326
rect 23945 37302 23946 37326
rect 23894 37274 23946 37302
rect 66 35677 118 35737
rect 66 35537 69 35677
rect 69 35537 115 35677
rect 115 35537 118 35677
rect 66 35477 118 35537
rect 23894 35712 23946 35740
rect 23894 35688 23899 35712
rect 23899 35688 23945 35712
rect 23945 35688 23946 35712
rect 23894 35502 23899 35522
rect 23899 35502 23945 35522
rect 23945 35502 23946 35522
rect 23894 35470 23946 35502
rect 66 33877 118 33937
rect 66 33737 69 33877
rect 69 33737 115 33877
rect 115 33737 118 33877
rect 66 33677 118 33737
rect 23894 33912 23946 33944
rect 23894 33892 23899 33912
rect 23899 33892 23945 33912
rect 23945 33892 23946 33912
rect 23894 33702 23899 33726
rect 23899 33702 23945 33726
rect 23945 33702 23946 33726
rect 23894 33674 23946 33702
rect 66 32077 118 32137
rect 66 31937 69 32077
rect 69 31937 115 32077
rect 115 31937 118 32077
rect 66 31877 118 31937
rect 23894 32112 23946 32140
rect 23894 32088 23899 32112
rect 23899 32088 23945 32112
rect 23945 32088 23946 32112
rect 23894 31902 23899 31922
rect 23899 31902 23945 31922
rect 23945 31902 23946 31922
rect 23894 31870 23946 31902
rect 23894 30555 23946 30607
rect 23894 30388 23946 30389
rect 23894 30342 23899 30388
rect 23899 30342 23945 30388
rect 23945 30342 23946 30388
rect 23894 30337 23946 30342
rect 948 29803 1104 29818
rect 11742 29803 11898 29818
rect 948 29766 1033 29803
rect 1033 29766 1079 29803
rect 1079 29766 1104 29803
rect 11742 29766 11877 29803
rect 11877 29766 11898 29803
rect 22869 29766 23025 29818
rect 23369 28924 23421 28962
rect 23369 28910 23415 28924
rect 23415 28910 23421 28924
rect 23369 28724 23421 28776
rect 23386 28359 23415 28372
rect 23415 28359 23438 28372
rect 23386 28224 23438 28359
rect 23386 28216 23415 28224
rect 23415 28216 23438 28224
rect 23347 27584 23369 27593
rect 23369 27584 23399 27593
rect 23347 27449 23399 27584
rect 23347 27437 23369 27449
rect 23369 27437 23399 27449
rect 23156 26249 23208 26405
rect 23580 26249 23632 26405
rect 23571 25201 23623 25357
rect 23349 23880 23369 23922
rect 23369 23880 23401 23922
rect 23349 23766 23401 23880
rect 23578 22170 23630 22222
rect 23764 22170 23816 22222
rect 23536 21972 23588 22024
rect 23156 21768 23208 21820
rect 23364 20127 23416 20179
rect 23314 19951 23470 19984
rect 23314 19932 23369 19951
rect 23369 19932 23415 19951
rect 23415 19932 23470 19951
rect 23139 18131 23191 18183
rect 23319 18174 23371 18183
rect 23319 18131 23363 18174
rect 23363 18131 23371 18174
rect 23295 17936 23347 17988
rect 23443 17719 23495 17823
rect 23443 17673 23472 17719
rect 23472 17673 23495 17719
rect 23443 17667 23495 17673
rect 23366 16923 23418 16939
rect 23366 16887 23418 16923
rect 23216 15608 23268 15609
rect 23216 15562 23222 15608
rect 23222 15562 23268 15608
rect 23216 15557 23268 15562
rect 23402 15557 23454 15609
rect 23164 15007 23168 15015
rect 23168 15007 23214 15015
rect 23214 15007 23216 15015
rect 23164 14963 23216 15007
rect 23164 14797 23168 14829
rect 23168 14797 23214 14829
rect 23214 14797 23216 14829
rect 23164 14777 23216 14797
rect 23612 15007 23616 15015
rect 23616 15007 23662 15015
rect 23662 15007 23664 15015
rect 23612 14963 23664 15007
rect 23612 14797 23616 14829
rect 23616 14797 23662 14829
rect 23662 14797 23664 14829
rect 23612 14777 23664 14797
rect 23169 12524 23221 12576
rect 23169 12338 23172 12390
rect 23172 12338 23218 12390
rect 23218 12338 23221 12390
rect 23169 11986 23172 12038
rect 23172 11986 23218 12038
rect 23218 11986 23221 12038
rect 23169 11800 23172 11852
rect 23172 11800 23218 11852
rect 23218 11800 23221 11852
rect 23395 12524 23447 12576
rect 23395 12306 23396 12358
rect 23396 12306 23442 12358
rect 23442 12306 23447 12358
rect 23395 12088 23396 12140
rect 23396 12088 23442 12140
rect 23442 12088 23447 12140
rect 23395 11871 23396 11923
rect 23396 11871 23442 11923
rect 23442 11871 23447 11923
rect 23610 12524 23662 12576
rect 23610 12338 23620 12390
rect 23620 12338 23662 12390
rect 23610 11986 23620 12038
rect 23620 11986 23662 12038
rect 23610 11800 23620 11852
rect 23620 11800 23662 11852
rect 23395 11653 23396 11705
rect 23396 11653 23442 11705
rect 23442 11653 23447 11705
rect 23169 11381 23172 11433
rect 23172 11381 23218 11433
rect 23218 11381 23221 11433
rect 23169 11195 23172 11247
rect 23172 11195 23218 11247
rect 23218 11195 23221 11247
rect 23395 11435 23396 11487
rect 23396 11435 23442 11487
rect 23442 11435 23447 11487
rect 23395 11218 23396 11270
rect 23396 11218 23442 11270
rect 23442 11218 23447 11270
rect 23610 11381 23620 11433
rect 23620 11381 23662 11433
rect 23610 11195 23620 11247
rect 23620 11195 23662 11247
rect 23395 11000 23396 11052
rect 23396 11000 23442 11052
rect 23442 11000 23447 11052
rect 23395 10817 23396 10835
rect 23396 10817 23442 10835
rect 23442 10817 23447 10835
rect 23395 10783 23447 10817
rect 23395 10565 23447 10617
rect 23395 10361 23396 10399
rect 23396 10361 23442 10399
rect 23442 10361 23447 10399
rect 23395 10347 23447 10361
rect 23395 10155 23396 10182
rect 23396 10155 23442 10182
rect 23442 10155 23447 10182
rect 23395 10130 23447 10155
rect 23395 9949 23396 9964
rect 23396 9949 23442 9964
rect 23442 9949 23447 9964
rect 23395 9912 23447 9949
rect 23395 9743 23396 9746
rect 23396 9743 23442 9746
rect 23442 9743 23447 9746
rect 23395 9694 23447 9743
rect 23395 9480 23447 9529
rect 23395 9477 23396 9480
rect 23396 9477 23442 9480
rect 23442 9477 23447 9480
rect 23395 9274 23447 9311
rect 23395 9259 23396 9274
rect 23396 9259 23442 9274
rect 23442 9259 23447 9274
rect 23395 9068 23447 9093
rect 23395 9041 23396 9068
rect 23396 9041 23442 9068
rect 23442 9041 23447 9068
rect 23395 8862 23447 8876
rect 23395 8824 23396 8862
rect 23396 8824 23442 8862
rect 23442 8824 23447 8862
rect 23395 8606 23396 8658
rect 23396 8606 23442 8658
rect 23442 8606 23447 8658
rect 23173 7722 23225 7774
rect 23173 7536 23225 7588
rect 23173 7350 23225 7402
rect 23395 8408 23396 8441
rect 23396 8408 23442 8441
rect 23442 8408 23447 8441
rect 23395 8389 23447 8408
rect 23395 8171 23447 8223
rect 23395 7953 23447 8005
rect 23395 7736 23447 7788
rect 23395 7518 23447 7570
rect 23395 7300 23447 7352
rect 23615 7722 23667 7774
rect 23615 7536 23667 7588
rect 23615 7350 23667 7402
rect 23297 4921 23349 4973
rect 23509 4921 23561 4973
rect 23297 4703 23349 4755
rect 23509 4703 23561 4755
<< metal2 >>
rect 54 89535 130 89547
rect 54 89275 66 89535
rect 118 89275 130 89535
rect 54 87936 130 89275
rect 54 87676 66 87936
rect 118 87676 130 87936
rect 54 86137 130 87676
rect 23857 89477 23982 89517
rect 23857 89425 23894 89477
rect 23946 89425 23982 89477
rect 23857 89259 23982 89425
rect 23857 89207 23894 89259
rect 23946 89207 23982 89259
rect 23857 87940 23982 89207
rect 23857 87888 23894 87940
rect 23946 87888 23982 87940
rect 23857 87722 23982 87888
rect 23857 87670 23894 87722
rect 23946 87670 23982 87722
rect 23857 87576 23982 87670
rect 54 85877 66 86137
rect 118 85877 130 86137
rect 54 84337 130 85877
rect 54 84077 66 84337
rect 118 84077 130 84337
rect 54 82537 130 84077
rect 54 82277 66 82537
rect 118 82277 130 82537
rect 54 80736 130 82277
rect 54 80476 66 80736
rect 118 80476 130 80736
rect 54 78937 130 80476
rect 54 78677 66 78937
rect 118 78677 130 78937
rect 54 77138 130 78677
rect 54 76878 66 77138
rect 118 76878 130 77138
rect 54 75337 130 76878
rect 54 75077 66 75337
rect 118 75077 130 75337
rect 54 73537 130 75077
rect 54 73277 66 73537
rect 118 73277 130 73537
rect 54 71737 130 73277
rect 54 71477 66 71737
rect 118 71477 130 71737
rect 54 69937 130 71477
rect 54 69677 66 69937
rect 118 69677 130 69937
rect 54 68137 130 69677
rect 54 67877 66 68137
rect 118 67877 130 68137
rect 54 66337 130 67877
rect 54 66077 66 66337
rect 118 66077 130 66337
rect 54 64537 130 66077
rect 54 64277 66 64537
rect 118 64277 130 64537
rect 54 62737 130 64277
rect 54 62477 66 62737
rect 118 62477 130 62737
rect 54 60937 130 62477
rect 54 60677 66 60937
rect 118 60677 130 60937
rect 54 59137 130 60677
rect 54 58877 66 59137
rect 118 58877 130 59137
rect 54 57337 130 58877
rect 54 57077 66 57337
rect 118 57077 130 57337
rect 54 55537 130 57077
rect 54 55277 66 55537
rect 118 55277 130 55537
rect 54 53749 130 55277
rect 50 53737 130 53749
rect 50 53477 62 53737
rect 114 53477 130 53737
rect 50 53465 130 53477
rect 54 51937 130 53465
rect 54 51677 66 51937
rect 118 51677 130 51937
rect 54 50137 130 51677
rect 54 49877 66 50137
rect 118 49877 130 50137
rect 54 48337 130 49877
rect 54 48077 66 48337
rect 118 48077 130 48337
rect 54 46537 130 48077
rect 54 46277 66 46537
rect 118 46277 130 46537
rect 54 44737 130 46277
rect 54 44477 66 44737
rect 118 44477 130 44737
rect 54 42937 130 44477
rect 54 42677 66 42937
rect 118 42677 130 42937
rect 54 41137 130 42677
rect 54 40877 66 41137
rect 118 40877 130 41137
rect 54 39337 130 40877
rect 54 39077 66 39337
rect 118 39077 130 39337
rect 54 37537 130 39077
rect 54 37277 66 37537
rect 118 37277 130 37537
rect 54 35737 130 37277
rect 54 35477 66 35737
rect 118 35477 130 35737
rect 54 33937 130 35477
rect 54 33677 66 33937
rect 118 33677 130 33937
rect 54 32137 130 33677
rect 54 31877 66 32137
rect 118 31877 130 32137
rect 54 30241 130 31877
rect 23857 86140 23982 86219
rect 23857 86088 23894 86140
rect 23946 86088 23982 86140
rect 23857 85922 23982 86088
rect 23857 85870 23894 85922
rect 23946 85870 23982 85922
rect 23857 84340 23982 85870
rect 23857 84288 23894 84340
rect 23946 84288 23982 84340
rect 23857 84122 23982 84288
rect 23857 84070 23894 84122
rect 23946 84070 23982 84122
rect 23857 82540 23982 84070
rect 23857 82488 23894 82540
rect 23946 82488 23982 82540
rect 23857 82322 23982 82488
rect 23857 82270 23894 82322
rect 23946 82270 23982 82322
rect 23857 80740 23982 82270
rect 23857 80688 23894 80740
rect 23946 80688 23982 80740
rect 23857 80522 23982 80688
rect 23857 80470 23894 80522
rect 23946 80470 23982 80522
rect 23857 78940 23982 80470
rect 23857 78888 23894 78940
rect 23946 78888 23982 78940
rect 23857 78722 23982 78888
rect 23857 78670 23894 78722
rect 23946 78670 23982 78722
rect 23857 77140 23982 78670
rect 23857 77088 23894 77140
rect 23946 77088 23982 77140
rect 23857 76922 23982 77088
rect 23857 76870 23894 76922
rect 23946 76870 23982 76922
rect 23857 75340 23982 76870
rect 23857 75288 23894 75340
rect 23946 75288 23982 75340
rect 23857 75122 23982 75288
rect 23857 75070 23894 75122
rect 23946 75070 23982 75122
rect 23857 73540 23982 75070
rect 23857 73488 23894 73540
rect 23946 73488 23982 73540
rect 23857 73322 23982 73488
rect 23857 73270 23894 73322
rect 23946 73270 23982 73322
rect 23857 71740 23982 73270
rect 23857 71688 23894 71740
rect 23946 71688 23982 71740
rect 23857 71522 23982 71688
rect 23857 71470 23894 71522
rect 23946 71470 23982 71522
rect 23857 69940 23982 71470
rect 23857 69888 23894 69940
rect 23946 69888 23982 69940
rect 23857 69722 23982 69888
rect 23857 69670 23894 69722
rect 23946 69670 23982 69722
rect 23857 68140 23982 69670
rect 23857 68088 23894 68140
rect 23946 68088 23982 68140
rect 23857 67922 23982 68088
rect 23857 67870 23894 67922
rect 23946 67870 23982 67922
rect 23857 66340 23982 67870
rect 23857 66288 23894 66340
rect 23946 66288 23982 66340
rect 23857 66122 23982 66288
rect 23857 66070 23894 66122
rect 23946 66070 23982 66122
rect 23857 64540 23982 66070
rect 23857 64488 23894 64540
rect 23946 64488 23982 64540
rect 23857 64322 23982 64488
rect 23857 64270 23894 64322
rect 23946 64270 23982 64322
rect 23857 62740 23982 64270
rect 23857 62688 23894 62740
rect 23946 62688 23982 62740
rect 23857 62522 23982 62688
rect 23857 62470 23894 62522
rect 23946 62470 23982 62522
rect 23857 60940 23982 62470
rect 23857 60888 23894 60940
rect 23946 60888 23982 60940
rect 23857 60722 23982 60888
rect 23857 60670 23894 60722
rect 23946 60670 23982 60722
rect 23857 59140 23982 60670
rect 23857 59088 23894 59140
rect 23946 59088 23982 59140
rect 23857 58922 23982 59088
rect 23857 58870 23894 58922
rect 23946 58870 23982 58922
rect 23857 57340 23982 58870
rect 23857 57288 23894 57340
rect 23946 57288 23982 57340
rect 23857 57122 23982 57288
rect 23857 57070 23894 57122
rect 23946 57070 23982 57122
rect 23857 55544 23982 57070
rect 23857 55492 23894 55544
rect 23946 55492 23982 55544
rect 23857 55326 23982 55492
rect 23857 55274 23894 55326
rect 23946 55274 23982 55326
rect 23857 53740 23982 55274
rect 23857 53688 23894 53740
rect 23946 53688 23982 53740
rect 23857 53522 23982 53688
rect 23857 53470 23894 53522
rect 23946 53470 23982 53522
rect 23857 51944 23982 53470
rect 23857 51892 23894 51944
rect 23946 51892 23982 51944
rect 23857 51726 23982 51892
rect 23857 51674 23894 51726
rect 23946 51674 23982 51726
rect 23857 50140 23982 51674
rect 23857 50088 23894 50140
rect 23946 50088 23982 50140
rect 23857 49922 23982 50088
rect 23857 49870 23894 49922
rect 23946 49870 23982 49922
rect 23857 48344 23982 49870
rect 23857 48292 23894 48344
rect 23946 48292 23982 48344
rect 23857 48126 23982 48292
rect 23857 48074 23894 48126
rect 23946 48074 23982 48126
rect 23857 46540 23982 48074
rect 23857 46488 23894 46540
rect 23946 46488 23982 46540
rect 23857 46322 23982 46488
rect 23857 46270 23894 46322
rect 23946 46270 23982 46322
rect 23857 44744 23982 46270
rect 23857 44692 23894 44744
rect 23946 44692 23982 44744
rect 23857 44526 23982 44692
rect 23857 44474 23894 44526
rect 23946 44474 23982 44526
rect 23857 42940 23982 44474
rect 23857 42888 23894 42940
rect 23946 42888 23982 42940
rect 23857 42722 23982 42888
rect 23857 42670 23894 42722
rect 23946 42670 23982 42722
rect 23857 41144 23982 42670
rect 23857 41092 23894 41144
rect 23946 41092 23982 41144
rect 23857 40926 23982 41092
rect 23857 40874 23894 40926
rect 23946 40874 23982 40926
rect 23857 39340 23982 40874
rect 23857 39288 23894 39340
rect 23946 39288 23982 39340
rect 23857 39122 23982 39288
rect 23857 39070 23894 39122
rect 23946 39070 23982 39122
rect 23857 37544 23982 39070
rect 23857 37492 23894 37544
rect 23946 37492 23982 37544
rect 23857 37326 23982 37492
rect 23857 37274 23894 37326
rect 23946 37274 23982 37326
rect 23857 35740 23982 37274
rect 23857 35688 23894 35740
rect 23946 35688 23982 35740
rect 23857 35522 23982 35688
rect 23857 35470 23894 35522
rect 23946 35470 23982 35522
rect 23857 33944 23982 35470
rect 23857 33892 23894 33944
rect 23946 33892 23982 33944
rect 23857 33726 23982 33892
rect 23857 33674 23894 33726
rect 23946 33674 23982 33726
rect 23857 32140 23982 33674
rect 23857 32088 23894 32140
rect 23946 32088 23982 32140
rect 23857 31922 23982 32088
rect 23857 31870 23894 31922
rect 23946 31870 23982 31922
rect -51 30231 233 30241
rect -51 30175 -41 30231
rect 223 30175 233 30231
rect -51 30165 233 30175
rect 977 29987 1077 31182
rect 977 29931 996 29987
rect 1052 29931 1077 29987
rect 977 29855 1077 29931
rect 977 29830 996 29855
rect 936 29818 996 29830
rect 1052 29830 1077 29855
rect 1052 29818 1116 29830
rect 936 29766 948 29818
rect 1104 29766 1116 29818
rect 936 29754 1116 29766
rect 977 29723 1077 29754
rect 977 29667 996 29723
rect 1052 29667 1077 29723
rect 977 29591 1077 29667
rect 977 29535 996 29591
rect 1052 29535 1077 29591
rect 977 29471 1077 29535
rect 1337 29071 1437 31182
rect 11777 29987 11877 31182
rect 11777 29931 11798 29987
rect 11854 29931 11877 29987
rect 11777 29855 11877 29931
rect 11777 29830 11798 29855
rect 11730 29818 11798 29830
rect 11854 29830 11877 29855
rect 11854 29818 11910 29830
rect 11730 29766 11742 29818
rect 11898 29766 11910 29818
rect 11730 29754 11910 29766
rect 11777 29723 11877 29754
rect 11777 29667 11798 29723
rect 11854 29667 11877 29723
rect 11777 29591 11877 29667
rect 11777 29535 11798 29591
rect 11854 29535 11877 29591
rect 11777 29517 11877 29535
rect 1337 29015 1358 29071
rect 1414 29015 1437 29071
rect 1337 28939 1437 29015
rect 1337 28883 1358 28939
rect 1414 28883 1437 28939
rect 1337 28807 1437 28883
rect 1337 28751 1358 28807
rect 1414 28751 1437 28807
rect 1337 28675 1437 28751
rect 1337 28619 1358 28675
rect 1414 28619 1437 28675
rect 1337 28543 1437 28619
rect 1337 28487 1358 28543
rect 1414 28487 1437 28543
rect 1337 28411 1437 28487
rect 1337 28355 1358 28411
rect 1414 28355 1437 28411
rect 1337 28279 1437 28355
rect 1337 28223 1358 28279
rect 1414 28223 1437 28279
rect 1337 28147 1437 28223
rect 1337 28091 1358 28147
rect 1414 28091 1437 28147
rect 1337 28015 1437 28091
rect 1337 27959 1358 28015
rect 1414 27959 1437 28015
rect 1337 27883 1437 27959
rect 1337 27827 1358 27883
rect 1414 27827 1437 27883
rect 1337 27751 1437 27827
rect 1337 27695 1358 27751
rect 1414 27695 1437 27751
rect 1337 27619 1437 27695
rect 1337 27563 1358 27619
rect 1414 27563 1437 27619
rect 1337 27527 1437 27563
rect 12137 29071 12237 31182
rect 12137 29015 12158 29071
rect 12214 29015 12237 29071
rect 12137 28939 12237 29015
rect 12137 28883 12158 28939
rect 12214 28883 12237 28939
rect 12137 28807 12237 28883
rect 12137 28751 12158 28807
rect 12214 28751 12237 28807
rect 12137 28675 12237 28751
rect 12137 28619 12158 28675
rect 12214 28619 12237 28675
rect 12137 28543 12237 28619
rect 12137 28487 12158 28543
rect 12214 28487 12237 28543
rect 12137 28411 12237 28487
rect 12137 28355 12158 28411
rect 12214 28355 12237 28411
rect 12137 28279 12237 28355
rect 12137 28223 12158 28279
rect 12214 28223 12237 28279
rect 12137 28147 12237 28223
rect 12137 28091 12158 28147
rect 12214 28091 12237 28147
rect 12137 28015 12237 28091
rect 12137 27959 12158 28015
rect 12214 27959 12237 28015
rect 12137 27883 12237 27959
rect 12137 27827 12158 27883
rect 12214 27827 12237 27883
rect 12137 27751 12237 27827
rect 12137 27695 12158 27751
rect 12214 27695 12237 27751
rect 12137 27619 12237 27695
rect 12137 27563 12158 27619
rect 12214 27563 12237 27619
rect 12137 27527 12237 27563
rect 22577 29071 22677 31182
rect 22937 29987 23037 31182
rect 23857 30607 23982 31870
rect 23857 30555 23894 30607
rect 23946 30555 23982 30607
rect 22937 29931 22958 29987
rect 23014 29931 23037 29987
rect 22937 29855 23037 29931
rect 22937 29830 22958 29855
rect 22857 29818 22958 29830
rect 23014 29818 23037 29855
rect 22857 29766 22869 29818
rect 23025 29766 23037 29818
rect 22857 29754 23037 29766
rect 22577 29015 22598 29071
rect 22654 29015 22677 29071
rect 22577 28939 22677 29015
rect 22577 28883 22598 28939
rect 22654 28883 22677 28939
rect 22577 28807 22677 28883
rect 22577 28751 22598 28807
rect 22654 28751 22677 28807
rect 22577 28675 22677 28751
rect 22577 28619 22598 28675
rect 22654 28619 22677 28675
rect 22577 28543 22677 28619
rect 22577 28487 22598 28543
rect 22654 28487 22677 28543
rect 22577 28411 22677 28487
rect 22577 28355 22598 28411
rect 22654 28355 22677 28411
rect 22577 28279 22677 28355
rect 22577 28223 22598 28279
rect 22654 28223 22677 28279
rect 22577 28147 22677 28223
rect 22577 28091 22598 28147
rect 22654 28091 22677 28147
rect 22577 28015 22677 28091
rect 22577 27959 22598 28015
rect 22654 27959 22677 28015
rect 22577 27883 22677 27959
rect 22577 27827 22598 27883
rect 22654 27827 22677 27883
rect 22577 27751 22677 27827
rect 22577 27695 22598 27751
rect 22654 27695 22677 27751
rect 22577 27619 22677 27695
rect 22577 27563 22598 27619
rect 22654 27563 22677 27619
rect 22577 27527 22677 27563
rect 22937 29723 23037 29754
rect 22937 29667 22958 29723
rect 23014 29667 23037 29723
rect 22937 29591 23037 29667
rect 22937 29535 22958 29591
rect 23014 29535 23037 29591
rect 22937 27527 23037 29535
rect 23197 29350 23317 30533
rect 23154 29252 23317 29350
rect 23497 29350 23617 30533
rect 23857 30389 23982 30555
rect 23857 30337 23894 30389
rect 23946 30337 23982 30389
rect 23857 30297 23982 30337
rect 23497 29252 23625 29350
rect 23154 27543 23210 29252
rect 23328 28964 23456 28986
rect 23328 28908 23367 28964
rect 23423 28908 23456 28964
rect 23328 28778 23456 28908
rect 23328 28722 23367 28778
rect 23423 28722 23456 28778
rect 23328 28703 23456 28722
rect 23374 28372 23450 28384
rect 23374 28216 23386 28372
rect 23438 28322 23450 28372
rect 23569 28322 23625 29252
rect 23438 28266 23625 28322
rect 23438 28216 23450 28266
rect 23374 28204 23450 28216
rect 23335 27593 23411 27605
rect 23335 27543 23347 27593
rect 23154 27487 23347 27543
rect 23154 26417 23210 27487
rect 23335 27437 23347 27487
rect 23399 27437 23411 27593
rect 23335 27425 23411 27437
rect 23569 26417 23625 28266
rect 23144 26405 23220 26417
rect 23144 26249 23156 26405
rect 23208 26249 23220 26405
rect 23144 26237 23220 26249
rect 23568 26405 23644 26417
rect 23568 26249 23580 26405
rect 23632 26249 23644 26405
rect 23568 26237 23644 26249
rect 23154 21832 23210 26237
rect 23569 25369 23625 26237
rect 23559 25357 23635 25369
rect 23559 25201 23571 25357
rect 23623 25201 23635 25357
rect 23559 25189 23635 25201
rect 23337 23922 23413 23934
rect 23337 23766 23349 23922
rect 23401 23766 23413 23922
rect 23337 23754 23413 23766
rect 23144 21820 23220 21832
rect 23144 21768 23156 21820
rect 23208 21768 23220 21820
rect 23144 21756 23220 21768
rect 23347 21571 23403 23754
rect 23569 22344 23625 25189
rect 23548 22222 23856 22242
rect 23548 22170 23578 22222
rect 23630 22170 23764 22222
rect 23816 22170 23856 22222
rect 23548 22150 23856 22170
rect 23497 22026 23626 22065
rect 23497 21970 23534 22026
rect 23590 21970 23626 22026
rect 23497 21931 23626 21970
rect 23498 21808 23626 21931
rect 23498 21752 23534 21808
rect 23590 21752 23626 21808
rect 23498 21714 23626 21752
rect 23347 21515 23621 21571
rect 23129 20179 23452 20203
rect 23129 20127 23364 20179
rect 23416 20127 23452 20179
rect 23129 20106 23452 20127
rect 23129 18612 23221 20106
rect 23565 19996 23621 21515
rect 23302 19984 23621 19996
rect 23302 19932 23314 19984
rect 23470 19932 23621 19984
rect 23302 19920 23621 19932
rect 23129 18515 23320 18612
rect 23227 18206 23320 18515
rect 23101 18185 23409 18206
rect 23101 18129 23137 18185
rect 23193 18129 23317 18185
rect 23373 18129 23409 18185
rect 23101 18109 23409 18129
rect 23227 18011 23320 18109
rect 23227 17988 23386 18011
rect 23227 17936 23295 17988
rect 23347 17936 23386 17988
rect 23227 17914 23386 17936
rect 23565 17835 23621 19920
rect 23431 17823 23621 17835
rect 23431 17667 23443 17823
rect 23495 17779 23621 17823
rect 23495 17667 23507 17779
rect 23431 17655 23507 17667
rect 23328 16941 23456 17037
rect 23328 16885 23364 16941
rect 23420 16885 23456 16941
rect 23328 16808 23456 16885
rect 23768 16758 23856 22150
rect 23186 15611 23494 15629
rect 23186 15555 23214 15611
rect 23270 15555 23400 15611
rect 23456 15555 23494 15611
rect 23186 15537 23494 15555
rect 23144 15017 23236 15045
rect 23144 14961 23162 15017
rect 23218 14961 23236 15017
rect 23144 14831 23236 14961
rect 23144 14775 23162 14831
rect 23218 14775 23236 14831
rect 23144 14737 23236 14775
rect 23592 15017 23684 15045
rect 23592 14961 23610 15017
rect 23666 14961 23684 15017
rect 23592 14831 23684 14961
rect 23592 14775 23610 14831
rect 23666 14775 23684 14831
rect 23592 14737 23684 14775
rect 23149 12578 23241 12606
rect 23149 12522 23167 12578
rect 23223 12522 23241 12578
rect 23149 12392 23241 12522
rect 23149 12336 23167 12392
rect 23223 12336 23241 12392
rect 23149 12298 23241 12336
rect 23356 12576 23486 12616
rect 23356 12524 23395 12576
rect 23447 12524 23486 12576
rect 23356 12358 23486 12524
rect 23356 12306 23395 12358
rect 23447 12306 23486 12358
rect 23356 12140 23486 12306
rect 23590 12578 23682 12606
rect 23590 12522 23608 12578
rect 23664 12522 23682 12578
rect 23590 12392 23682 12522
rect 23590 12336 23608 12392
rect 23664 12336 23682 12392
rect 23590 12298 23682 12336
rect 23356 12088 23395 12140
rect 23447 12088 23486 12140
rect 23149 12040 23241 12068
rect 23149 11984 23167 12040
rect 23223 11984 23241 12040
rect 23149 11854 23241 11984
rect 23149 11798 23167 11854
rect 23223 11798 23241 11854
rect 23149 11760 23241 11798
rect 23356 11923 23486 12088
rect 23356 11871 23395 11923
rect 23447 11871 23486 11923
rect 23356 11705 23486 11871
rect 23590 12040 23682 12068
rect 23590 11984 23608 12040
rect 23664 11984 23682 12040
rect 23590 11854 23682 11984
rect 23590 11798 23608 11854
rect 23664 11798 23682 11854
rect 23590 11760 23682 11798
rect 23356 11653 23395 11705
rect 23447 11653 23486 11705
rect 23356 11487 23486 11653
rect 23149 11435 23241 11463
rect 23149 11379 23167 11435
rect 23223 11379 23241 11435
rect 23149 11249 23241 11379
rect 23149 11193 23167 11249
rect 23223 11193 23241 11249
rect 23149 11155 23241 11193
rect 23356 11435 23395 11487
rect 23447 11435 23486 11487
rect 23356 11270 23486 11435
rect 23356 11218 23395 11270
rect 23447 11218 23486 11270
rect 23356 11052 23486 11218
rect 23590 11435 23682 11463
rect 23590 11379 23608 11435
rect 23664 11379 23682 11435
rect 23590 11249 23682 11379
rect 23590 11193 23608 11249
rect 23664 11193 23682 11249
rect 23590 11155 23682 11193
rect 23356 11000 23395 11052
rect 23447 11000 23486 11052
rect 23356 10835 23486 11000
rect 23356 10783 23395 10835
rect 23447 10783 23486 10835
rect 23356 10617 23486 10783
rect 23356 10565 23395 10617
rect 23447 10565 23486 10617
rect 23356 10399 23486 10565
rect 23356 10347 23395 10399
rect 23447 10347 23486 10399
rect 23356 10182 23486 10347
rect 23356 10130 23395 10182
rect 23447 10130 23486 10182
rect 23356 9964 23486 10130
rect 23356 9912 23395 9964
rect 23447 9912 23486 9964
rect 23356 9746 23486 9912
rect 23356 9694 23395 9746
rect 23447 9694 23486 9746
rect 23356 9529 23486 9694
rect 23356 9477 23395 9529
rect 23447 9477 23486 9529
rect 23356 9311 23486 9477
rect 23356 9259 23395 9311
rect 23447 9259 23486 9311
rect 23356 9093 23486 9259
rect 23356 9041 23395 9093
rect 23447 9041 23486 9093
rect 23356 8876 23486 9041
rect 23356 8824 23395 8876
rect 23447 8824 23486 8876
rect 23356 8658 23486 8824
rect 23356 8606 23395 8658
rect 23447 8606 23486 8658
rect 23356 8441 23486 8606
rect 23356 8389 23395 8441
rect 23447 8389 23486 8441
rect 23356 8223 23486 8389
rect 23356 8171 23395 8223
rect 23447 8171 23486 8223
rect 23356 8005 23486 8171
rect 23356 7953 23395 8005
rect 23447 7953 23486 8005
rect 23153 7776 23245 7804
rect 23153 7720 23171 7776
rect 23227 7720 23245 7776
rect 23153 7590 23245 7720
rect 23153 7534 23171 7590
rect 23227 7534 23245 7590
rect 23153 7404 23245 7534
rect 23153 7348 23171 7404
rect 23227 7348 23245 7404
rect 23153 7310 23245 7348
rect 23356 7788 23486 7953
rect 23356 7736 23395 7788
rect 23447 7736 23486 7788
rect 23356 7570 23486 7736
rect 23356 7518 23395 7570
rect 23447 7518 23486 7570
rect 23356 7352 23486 7518
rect 23356 7300 23395 7352
rect 23447 7300 23486 7352
rect 23595 7776 23687 7804
rect 23595 7720 23613 7776
rect 23669 7720 23687 7776
rect 23595 7590 23687 7720
rect 23595 7534 23613 7590
rect 23669 7534 23687 7590
rect 23595 7404 23687 7534
rect 23595 7348 23613 7404
rect 23669 7348 23687 7404
rect 23595 7310 23687 7348
rect 23356 5014 23486 7300
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4757 23599 4919
rect 23259 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 23259 4662 23599 4701
<< via2 >>
rect -41 30175 223 30231
rect 996 29931 1052 29987
rect 996 29818 1052 29855
rect 996 29799 1052 29818
rect 996 29667 1052 29723
rect 996 29535 1052 29591
rect 11798 29931 11854 29987
rect 11798 29818 11854 29855
rect 11798 29799 11854 29818
rect 11798 29667 11854 29723
rect 11798 29535 11854 29591
rect 1358 29015 1414 29071
rect 1358 28883 1414 28939
rect 1358 28751 1414 28807
rect 1358 28619 1414 28675
rect 1358 28487 1414 28543
rect 1358 28355 1414 28411
rect 1358 28223 1414 28279
rect 1358 28091 1414 28147
rect 1358 27959 1414 28015
rect 1358 27827 1414 27883
rect 1358 27695 1414 27751
rect 1358 27563 1414 27619
rect 12158 29015 12214 29071
rect 12158 28883 12214 28939
rect 12158 28751 12214 28807
rect 12158 28619 12214 28675
rect 12158 28487 12214 28543
rect 12158 28355 12214 28411
rect 12158 28223 12214 28279
rect 12158 28091 12214 28147
rect 12158 27959 12214 28015
rect 12158 27827 12214 27883
rect 12158 27695 12214 27751
rect 12158 27563 12214 27619
rect 22958 29931 23014 29987
rect 22958 29818 23014 29855
rect 22958 29799 23014 29818
rect 22598 29015 22654 29071
rect 22598 28883 22654 28939
rect 22598 28751 22654 28807
rect 22598 28619 22654 28675
rect 22598 28487 22654 28543
rect 22598 28355 22654 28411
rect 22598 28223 22654 28279
rect 22598 28091 22654 28147
rect 22598 27959 22654 28015
rect 22598 27827 22654 27883
rect 22598 27695 22654 27751
rect 22598 27563 22654 27619
rect 22958 29667 23014 29723
rect 22958 29535 23014 29591
rect 23367 28962 23423 28964
rect 23367 28910 23369 28962
rect 23369 28910 23421 28962
rect 23421 28910 23423 28962
rect 23367 28908 23423 28910
rect 23367 28776 23423 28778
rect 23367 28724 23369 28776
rect 23369 28724 23421 28776
rect 23421 28724 23423 28776
rect 23367 28722 23423 28724
rect 23534 22024 23590 22026
rect 23534 21972 23536 22024
rect 23536 21972 23588 22024
rect 23588 21972 23590 22024
rect 23534 21970 23590 21972
rect 23534 21752 23590 21808
rect 23137 18183 23193 18185
rect 23137 18131 23139 18183
rect 23139 18131 23191 18183
rect 23191 18131 23193 18183
rect 23137 18129 23193 18131
rect 23317 18183 23373 18185
rect 23317 18131 23319 18183
rect 23319 18131 23371 18183
rect 23371 18131 23373 18183
rect 23317 18129 23373 18131
rect 23364 16939 23420 16941
rect 23364 16887 23366 16939
rect 23366 16887 23418 16939
rect 23418 16887 23420 16939
rect 23364 16885 23420 16887
rect 23214 15609 23270 15611
rect 23214 15557 23216 15609
rect 23216 15557 23268 15609
rect 23268 15557 23270 15609
rect 23214 15555 23270 15557
rect 23400 15609 23456 15611
rect 23400 15557 23402 15609
rect 23402 15557 23454 15609
rect 23454 15557 23456 15609
rect 23400 15555 23456 15557
rect 23162 15015 23218 15017
rect 23162 14963 23164 15015
rect 23164 14963 23216 15015
rect 23216 14963 23218 15015
rect 23162 14961 23218 14963
rect 23162 14829 23218 14831
rect 23162 14777 23164 14829
rect 23164 14777 23216 14829
rect 23216 14777 23218 14829
rect 23162 14775 23218 14777
rect 23610 15015 23666 15017
rect 23610 14963 23612 15015
rect 23612 14963 23664 15015
rect 23664 14963 23666 15015
rect 23610 14961 23666 14963
rect 23610 14829 23666 14831
rect 23610 14777 23612 14829
rect 23612 14777 23664 14829
rect 23664 14777 23666 14829
rect 23610 14775 23666 14777
rect 23167 12576 23223 12578
rect 23167 12524 23169 12576
rect 23169 12524 23221 12576
rect 23221 12524 23223 12576
rect 23167 12522 23223 12524
rect 23167 12390 23223 12392
rect 23167 12338 23169 12390
rect 23169 12338 23221 12390
rect 23221 12338 23223 12390
rect 23167 12336 23223 12338
rect 23608 12576 23664 12578
rect 23608 12524 23610 12576
rect 23610 12524 23662 12576
rect 23662 12524 23664 12576
rect 23608 12522 23664 12524
rect 23608 12390 23664 12392
rect 23608 12338 23610 12390
rect 23610 12338 23662 12390
rect 23662 12338 23664 12390
rect 23608 12336 23664 12338
rect 23167 12038 23223 12040
rect 23167 11986 23169 12038
rect 23169 11986 23221 12038
rect 23221 11986 23223 12038
rect 23167 11984 23223 11986
rect 23167 11852 23223 11854
rect 23167 11800 23169 11852
rect 23169 11800 23221 11852
rect 23221 11800 23223 11852
rect 23167 11798 23223 11800
rect 23608 12038 23664 12040
rect 23608 11986 23610 12038
rect 23610 11986 23662 12038
rect 23662 11986 23664 12038
rect 23608 11984 23664 11986
rect 23608 11852 23664 11854
rect 23608 11800 23610 11852
rect 23610 11800 23662 11852
rect 23662 11800 23664 11852
rect 23608 11798 23664 11800
rect 23167 11433 23223 11435
rect 23167 11381 23169 11433
rect 23169 11381 23221 11433
rect 23221 11381 23223 11433
rect 23167 11379 23223 11381
rect 23167 11247 23223 11249
rect 23167 11195 23169 11247
rect 23169 11195 23221 11247
rect 23221 11195 23223 11247
rect 23167 11193 23223 11195
rect 23608 11433 23664 11435
rect 23608 11381 23610 11433
rect 23610 11381 23662 11433
rect 23662 11381 23664 11433
rect 23608 11379 23664 11381
rect 23608 11247 23664 11249
rect 23608 11195 23610 11247
rect 23610 11195 23662 11247
rect 23662 11195 23664 11247
rect 23608 11193 23664 11195
rect 23171 7774 23227 7776
rect 23171 7722 23173 7774
rect 23173 7722 23225 7774
rect 23225 7722 23227 7774
rect 23171 7720 23227 7722
rect 23171 7588 23227 7590
rect 23171 7536 23173 7588
rect 23173 7536 23225 7588
rect 23225 7536 23227 7588
rect 23171 7534 23227 7536
rect 23171 7402 23227 7404
rect 23171 7350 23173 7402
rect 23173 7350 23225 7402
rect 23225 7350 23227 7402
rect 23171 7348 23227 7350
rect 23613 7774 23669 7776
rect 23613 7722 23615 7774
rect 23615 7722 23667 7774
rect 23667 7722 23669 7774
rect 23613 7720 23669 7722
rect 23613 7588 23669 7590
rect 23613 7536 23615 7588
rect 23615 7536 23667 7588
rect 23667 7536 23669 7588
rect 23613 7534 23669 7536
rect 23613 7402 23669 7404
rect 23613 7350 23615 7402
rect 23615 7350 23667 7402
rect 23667 7350 23669 7402
rect 23613 7348 23669 7350
rect 23295 4973 23351 4975
rect 23295 4921 23297 4973
rect 23297 4921 23349 4973
rect 23349 4921 23351 4973
rect 23295 4919 23351 4921
rect 23507 4973 23563 4975
rect 23507 4921 23509 4973
rect 23509 4921 23561 4973
rect 23561 4921 23563 4973
rect 23507 4919 23563 4921
rect 23295 4755 23351 4757
rect 23295 4703 23297 4755
rect 23297 4703 23349 4755
rect 23349 4703 23351 4755
rect 23295 4701 23351 4703
rect 23507 4755 23563 4757
rect 23507 4703 23509 4755
rect 23509 4703 23561 4755
rect 23561 4703 23563 4755
rect 23507 4701 23563 4703
<< metal3 >>
rect -1 89507 23681 89707
rect -1 30537 23681 30897
rect -51 30231 23681 30279
rect -51 30175 -41 30231
rect 223 30175 23681 30231
rect -51 30139 23681 30175
rect -1 29987 24087 29997
rect -1 29931 996 29987
rect 1052 29931 11798 29987
rect 11854 29931 22958 29987
rect 23014 29931 24087 29987
rect -1 29855 24087 29931
rect -1 29799 996 29855
rect 1052 29799 11798 29855
rect 11854 29799 22958 29855
rect 23014 29799 24087 29855
rect -1 29723 24087 29799
rect -1 29667 996 29723
rect 1052 29667 11798 29723
rect 11854 29667 22958 29723
rect 23014 29667 24087 29723
rect -1 29591 24087 29667
rect -1 29535 996 29591
rect 1052 29535 11798 29591
rect 11854 29535 22958 29591
rect 23014 29535 24087 29591
rect -1 29517 24087 29535
rect 22636 29105 24206 29106
rect 800 29071 24206 29105
rect 800 29015 1358 29071
rect 1414 29015 12158 29071
rect 12214 29015 22598 29071
rect 22654 29015 24206 29071
rect 800 28964 24206 29015
rect 800 28939 23367 28964
rect 800 28883 1358 28939
rect 1414 28883 12158 28939
rect 12214 28883 22598 28939
rect 22654 28908 23367 28939
rect 23423 28908 24206 28964
rect 22654 28883 24206 28908
rect 800 28807 24206 28883
rect 800 28751 1358 28807
rect 1414 28751 12158 28807
rect 12214 28751 22598 28807
rect 22654 28778 24206 28807
rect 22654 28751 23367 28778
rect 800 28722 23367 28751
rect 23423 28722 24206 28778
rect 800 28675 24206 28722
rect 800 28619 1358 28675
rect 1414 28619 12158 28675
rect 12214 28619 22598 28675
rect 22654 28619 24206 28675
rect 800 28543 24206 28619
rect 800 28487 1358 28543
rect 1414 28487 12158 28543
rect 12214 28487 22598 28543
rect 22654 28487 24206 28543
rect 800 28411 24206 28487
rect 800 28355 1358 28411
rect 1414 28355 12158 28411
rect 12214 28355 22598 28411
rect 22654 28355 24206 28411
rect 800 28279 24206 28355
rect 800 28223 1358 28279
rect 1414 28223 12158 28279
rect 12214 28223 22598 28279
rect 22654 28223 24206 28279
rect 800 28147 24206 28223
rect 800 28091 1358 28147
rect 1414 28091 12158 28147
rect 12214 28091 22598 28147
rect 22654 28091 24206 28147
rect 800 28015 24206 28091
rect 800 27959 1358 28015
rect 1414 27959 12158 28015
rect 12214 27959 22598 28015
rect 22654 27959 24206 28015
rect 800 27883 24206 27959
rect 800 27827 1358 27883
rect 1414 27827 12158 27883
rect 12214 27827 22598 27883
rect 22654 27827 24206 27883
rect 800 27751 24206 27827
rect 800 27695 1358 27751
rect 1414 27695 12158 27751
rect 12214 27695 22598 27751
rect 22654 27695 24206 27751
rect 800 27619 24206 27695
rect 800 27563 1358 27619
rect 1414 27563 12158 27619
rect 12214 27563 22598 27619
rect 22654 27563 24206 27619
rect 800 27297 24206 27563
rect 800 27296 24087 27297
rect 22691 22026 24206 23393
rect 22691 21970 23534 22026
rect 23590 21970 24206 22026
rect 22691 21808 24206 21970
rect 22691 21752 23534 21808
rect 23590 21752 24206 21808
rect 22691 21416 24206 21752
rect 22586 21304 24206 21305
rect 1314 21090 24206 21304
rect 1314 21089 23252 21090
rect 22586 20983 24206 20984
rect 1314 20768 24206 20983
rect 1314 20767 23252 20768
rect 22586 20661 24206 20662
rect 1314 20447 24206 20661
rect 1314 20446 23252 20447
rect 22586 20339 24206 20340
rect 1314 20125 24206 20339
rect 1314 20124 23252 20125
rect 1314 19433 23889 19648
rect 1314 19432 23252 19433
rect 1314 19111 23889 19326
rect 1314 19110 23252 19111
rect 1314 18789 23889 19004
rect 22586 18682 23889 18683
rect 1314 18467 23889 18682
rect 1314 18185 23889 18361
rect 1314 18129 23137 18185
rect 23193 18129 23317 18185
rect 23373 18129 23889 18185
rect 1314 17919 23889 18129
rect 1314 17918 23252 17919
rect 1314 16941 24206 17263
rect 1314 16885 23364 16941
rect 23420 16885 24206 16941
rect 1314 16808 24206 16885
rect 1314 16807 23252 16808
rect 1314 15611 23710 15720
rect 1314 15555 23214 15611
rect 23270 15555 23400 15611
rect 23456 15555 23710 15611
rect 1314 15017 23710 15555
rect 1314 14961 23162 15017
rect 23218 14961 23610 15017
rect 23666 14961 23710 15017
rect 1314 14831 23710 14961
rect 1314 14775 23162 14831
rect 23218 14775 23610 14831
rect 23666 14775 23710 14831
rect 1314 12997 23710 14775
rect 1314 12996 23252 12997
rect 1314 12578 23710 12711
rect 1314 12522 23167 12578
rect 23223 12522 23608 12578
rect 23664 12522 23710 12578
rect 1314 12392 23710 12522
rect 1314 12336 23167 12392
rect 23223 12336 23608 12392
rect 23664 12336 23710 12392
rect 1314 12040 23710 12336
rect 1314 11984 23167 12040
rect 23223 11984 23608 12040
rect 23664 11984 23710 12040
rect 1314 11854 23710 11984
rect 1314 11798 23167 11854
rect 23223 11798 23608 11854
rect 23664 11798 23710 11854
rect 1314 11435 23710 11798
rect 1314 11379 23167 11435
rect 23223 11379 23608 11435
rect 23664 11379 23710 11435
rect 1314 11249 23710 11379
rect 1314 11193 23167 11249
rect 23223 11193 23608 11249
rect 23664 11193 23710 11249
rect 1314 9309 23710 11193
rect 1314 9308 23252 9309
rect 22658 9158 23710 9160
rect 1262 8442 23710 9158
rect 22658 7827 23710 7828
rect 1262 7776 24488 7827
rect 1262 7720 23171 7776
rect 23227 7720 23613 7776
rect 23669 7720 24488 7776
rect 1262 7590 24488 7720
rect 1262 7534 23171 7590
rect 23227 7534 23613 7590
rect 23669 7534 24488 7590
rect 1262 7404 24488 7534
rect 1262 7348 23171 7404
rect 23227 7348 23613 7404
rect 23669 7348 24488 7404
rect 1262 7016 24488 7348
rect 1314 5154 23971 6474
rect 1165 4923 22567 5011
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4758 23599 4919
rect 1165 4757 23599 4758
rect 1165 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 1165 4662 23599 4701
rect 1314 3133 24166 4495
rect 1314 1961 24276 2576
rect 1314 1286 23252 1855
rect 1314 747 24089 1179
rect 1314 155 24508 610
rect 1277 -959 24602 -504
rect 1277 -1599 23252 -1247
rect 1277 -2041 23252 -1953
rect 1277 -2517 23252 -2165
rect 1277 -3242 23252 -2787
use dcap_103_novia_512x8m81  dcap_103_novia_512x8m81_0
array 0 35 619 0 0 0
timestamp 1750858719
transform 1 0 288 0 1 29009
box 0 0 1 1
use M2_M1$$43374636_512x8m81  M2_M1$$43374636_512x8m81_0
timestamp 1750858719
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1750858719
transform -1 0 22947 0 -1 29792
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1750858719
transform -1 0 11820 0 -1 29792
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1750858719
transform -1 0 1026 0 -1 29792
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_0
timestamp 1750858719
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_0
timestamp 1750858719
transform 1 0 12186 0 1 28317
box 0 0 1 1
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_1
timestamp 1750858719
transform 1 0 22626 0 1 28317
box 0 0 1 1
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_2
timestamp 1750858719
transform 1 0 1386 0 1 28317
box 0 0 1 1
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_0
timestamp 1750858719
transform 1 0 1024 0 1 29761
box 0 0 1 1
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_1
timestamp 1750858719
transform 1 0 11826 0 1 29761
box 0 0 1 1
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_2
timestamp 1750858719
transform 1 0 22986 0 1 29761
box 0 0 1 1
use rarray4_512_512x8m81  rarray4_512_512x8m81_0
timestamp 1750858719
transform 1 0 907 0 1 31107
box -1997 -68 22836 57668
use rdummy_512x4_512x8m81  rdummy_512x4_512x8m81_0
timestamp 1750858719
transform 1 0 307 0 1 30207
box -219 -22942 23616 59468
use saout_m2_512x8m81  saout_m2_512x8m81_0
timestamp 1750858719
transform 1 0 11820 0 1 -1
box -269 -3393 7633 31140
use saout_m2_512x8m81  saout_m2_512x8m81_1
timestamp 1750858719
transform 1 0 1020 0 1 -1
box -269 -3393 7633 31140
use saout_R_m2_512x8m81  saout_R_m2_512x8m81_0
timestamp 1750858719
transform -1 0 12194 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_512x8m81  saout_R_m2_512x8m81_1
timestamp 1750858719
transform -1 0 22994 0 1 6
box -269 -3400 7633 31133
<< labels >>
rlabel metal3 s 1592 60366 1592 60366 4 WL[32]
port 1 nsew
rlabel metal3 s 1592 61266 1592 61266 4 WL[33]
port 2 nsew
rlabel metal3 s 1592 62166 1592 62166 4 WL[34]
port 3 nsew
rlabel metal3 s 1592 63066 1592 63066 4 WL[35]
port 4 nsew
rlabel metal3 s 1592 63966 1592 63966 4 WL[36]
port 5 nsew
rlabel metal3 s 1592 64866 1592 64866 4 WL[37]
port 6 nsew
rlabel metal3 s 1592 69366 1592 69366 4 WL[42]
port 7 nsew
rlabel metal3 s 1592 71166 1592 71166 4 WL[44]
port 8 nsew
rlabel metal3 s 1592 72966 1592 72966 4 WL[46]
port 9 nsew
rlabel metal3 s 1592 74766 1592 74766 4 WL[48]
port 10 nsew
rlabel metal3 s 1592 76566 1592 76566 4 WL[50]
port 11 nsew
rlabel metal3 s 1592 78366 1592 78366 4 WL[52]
port 12 nsew
rlabel metal3 s 1592 80166 1592 80166 4 WL[54]
port 13 nsew
rlabel metal3 s 1592 81966 1592 81966 4 WL[56]
port 14 nsew
rlabel metal3 s 1592 82866 1592 82866 4 WL[57]
port 15 nsew
rlabel metal3 s 1592 84666 1592 84666 4 WL[59]
port 16 nsew
rlabel metal3 s 1592 89157 1592 89157 4 DWL
port 17 nsew
rlabel metal3 s 1777 89717 1777 89717 4 VSS
port 18 nsew
rlabel metal3 s 1592 86465 1592 86465 4 WL[61]
port 19 nsew
rlabel metal3 s 1592 77465 1592 77465 4 WL[51]
port 20 nsew
rlabel metal3 s 1608 57668 1608 57668 4 WL[29]
port 21 nsew
rlabel metal3 s 1608 54068 1608 54068 4 WL[25]
port 22 nsew
rlabel metal3 s 1608 53168 1608 53168 4 WL[24]
port 23 nsew
rlabel metal3 s 1608 52268 1608 52268 4 WL[23]
port 24 nsew
rlabel metal3 s 1608 51368 1608 51368 4 WL[22]
port 25 nsew
rlabel metal3 s 1608 49568 1608 49568 4 WL[20]
port 26 nsew
rlabel metal3 s 1608 55868 1608 55868 4 WL[27]
port 27 nsew
rlabel metal3 s 1608 58568 1608 58568 4 WL[30]
port 28 nsew
rlabel metal3 s 1608 47768 1608 47768 4 WL[18]
port 29 nsew
rlabel metal3 s 1592 68465 1592 68465 4 WL[41]
port 30 nsew
rlabel metal3 s 1608 45068 1608 45068 4 WL[15]
port 31 nsew
rlabel metal3 s 1592 65765 1592 65765 4 WL[38]
port 32 nsew
rlabel metal3 s 1592 72065 1592 72065 4 WL[45]
port 33 nsew
rlabel metal3 s 1592 70265 1592 70265 4 WL[43]
port 34 nsew
rlabel metal3 s 1592 67565 1592 67565 4 WL[40]
port 35 nsew
rlabel metal3 s 1592 66665 1592 66665 4 WL[39]
port 36 nsew
rlabel metal3 s 1608 59468 1608 59468 4 WL[31]
port 37 nsew
rlabel metal3 s 1608 44168 1608 44168 4 WL[14]
port 38 nsew
rlabel metal3 s 1608 45968 1608 45968 4 WL[16]
port 39 nsew
rlabel metal3 s 1608 46868 1608 46868 4 WL[17]
port 40 nsew
rlabel metal3 s 1608 54968 1608 54968 4 WL[26]
port 41 nsew
rlabel metal3 s 1608 48668 1608 48668 4 WL[19]
port 42 nsew
rlabel metal3 s 1592 83765 1592 83765 4 WL[58]
port 43 nsew
rlabel metal3 s 1592 85565 1592 85565 4 WL[60]
port 44 nsew
rlabel metal3 s 1592 87365 1592 87365 4 WL[62]
port 45 nsew
rlabel metal3 s 1608 56768 1608 56768 4 WL[28]
port 46 nsew
rlabel metal3 s 1592 88265 1592 88265 4 WL[63]
port 47 nsew
rlabel metal3 s 1608 50468 1608 50468 4 WL[21]
port 48 nsew
rlabel metal3 s 1592 75665 1592 75665 4 WL[49]
port 49 nsew
rlabel metal3 s 1592 79265 1592 79265 4 WL[53]
port 50 nsew
rlabel metal3 s 1592 73865 1592 73865 4 WL[47]
port 51 nsew
rlabel metal3 s 1592 81065 1592 81065 4 WL[55]
port 52 nsew
rlabel metal3 s 240 30277 240 30277 4 VSS
port 18 nsew
rlabel metal3 s 1777 5806 1777 5806 4 VSS
port 18 nsew
rlabel metal3 s 1608 31568 1608 31568 4 WL[0]
port 53 nsew
rlabel metal3 s 1608 33368 1608 33368 4 WL[2]
port 54 nsew
rlabel metal3 s 1608 42368 1608 42368 4 WL[12]
port 55 nsew
rlabel metal3 s 1608 34268 1608 34268 4 WL[3]
port 56 nsew
rlabel metal3 s 1608 35168 1608 35168 4 WL[4]
port 57 nsew
flabel metal3 s 1659 -781 1659 -781 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
rlabel metal3 s 1608 37868 1608 37868 4 WL[7]
port 59 nsew
rlabel metal3 s 1608 38768 1608 38768 4 WL[8]
port 60 nsew
rlabel metal3 s 1608 39668 1608 39668 4 WL[9]
port 61 nsew
rlabel metal3 s 1608 32468 1608 32468 4 WL[1]
port 62 nsew
rlabel metal3 s 1705 21162 1705 21162 4 ypass[7]
port 63 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 64 nsew
flabel metal3 s 1659 -2347 1659 -2347 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 64 nsew
rlabel metal3 s 1607 36068 1607 36068 4 WL[5]
port 65 nsew
flabel metal3 s 1659 -1446 1659 -1446 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
rlabel metal3 s 1777 1467 1777 1467 4 men
port 64 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 64 nsew
rlabel metal3 s 1704 18591 1704 18591 4 ypass[0]
port 66 nsew
rlabel metal3 s 1608 40568 1608 40568 4 WL[10]
port 67 nsew
rlabel metal3 s 1608 43268 1608 43268 4 WL[13]
port 68 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 64 nsew
rlabel metal3 s 1704 18914 1704 18914 4 ypass[1]
port 69 nsew
rlabel metal3 s 1704 19231 1704 19231 4 ypass[2]
port 70 nsew
rlabel metal3 s 1704 19548 1704 19548 4 ypass[3]
port 71 nsew
rlabel metal3 s 1704 20204 1704 20204 4 ypass[4]
port 72 nsew
rlabel metal3 s 1704 20528 1704 20528 4 ypass[5]
port 73 nsew
rlabel metal3 s 1704 20845 1704 20845 4 ypass[6]
port 74 nsew
rlabel metal3 s 1774 1467 1774 1467 4 men
port 64 nsew
rlabel metal3 s 1607 36968 1607 36968 4 WL[6]
port 75 nsew
rlabel metal3 s 1346 4726 1346 4726 4 tblhl
port 76 nsew
flabel metal3 s 1659 -2004 1659 -2004 0 FreeSans 1000 0 0 0 GWEN
port 77 nsew
flabel metal3 s 1659 -3019 1659 -3019 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
rlabel metal3 s 1346 4983 1346 4983 4 GWE
port 78 nsew
rlabel metal3 s 1777 8832 1777 8832 4 VDD
port 58 nsew
rlabel metal3 s 1608 41468 1608 41468 4 WL[11]
port 79 nsew
flabel metal3 s 1659 390 1659 390 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 3623 1659 3623 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 7598 1659 7598 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 14001 1659 14001 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 18106 1659 18106 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 28191 1659 28191 0 FreeSans 1600 0 0 0 VDD
port 58 nsew
flabel metal3 s 315 29753 315 29753 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 23123 1659 23123 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 16976 1659 16976 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 12236 1659 12236 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 6155 1659 6155 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 2247 1659 2247 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 949 1659 949 0 FreeSans 1600 0 0 0 VSS
port 18 nsew
rlabel metal2 s 1525 104 1525 104 4 din[4]
port 80 nsew
rlabel metal2 s 22492 104 22492 104 4 din[7]
port 81 nsew
rlabel metal2 s 10847 138 10847 138 4 q[5]
port 82 nsew
rlabel metal2 s 13174 104 13174 104 4 q[6]
port 83 nsew
rlabel metal2 s 21634 104 21634 104 4 q[7]
port 84 nsew
rlabel metal2 s 11686 104 11686 104 4 din[5]
port 85 nsew
rlabel metal2 s 12325 104 12325 104 4 din[6]
port 86 nsew
rlabel metal2 s 2371 104 2371 104 4 q[4]
port 87 nsew
rlabel metal1 s 7342 15928 7342 15928 4 pcb[6]
port 88 nsew
rlabel metal1 s 5921 15928 5921 15928 4 pcb[7]
port 89 nsew
rlabel metal1 s 18209 15928 18209 15928 4 pcb[4]
port 90 nsew
rlabel metal1 s 1827 18163 1827 18163 4 vdd
port 91 nsew
flabel metal1 s 22465 -3332 22465 -3332 0 FreeSans 600 0 0 0 WEN[4]
port 92 nsew
flabel metal1 s 1584 -3332 1584 -3332 0 FreeSans 600 0 0 0 WEN[7]
port 93 nsew
rlabel metal1 s 16588 15928 16588 15928 4 pcb[5]
port 94 nsew
flabel metal1 s 12358 -3332 12358 -3332 0 FreeSans 600 0 0 0 WEN[5]
port 95 nsew
flabel metal1 s 11643 -3332 11643 -3332 0 FreeSans 600 0 0 0 WEN[6]
port 96 nsew
<< properties >>
string GDS_END 2831526
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2819152
<< end >>
