magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 1240 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 470 210 530 380
rect 700 210 760 380
rect 810 210 870 380
rect 980 210 1040 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 470 1110 530 1450
rect 700 1110 760 1450
rect 810 1110 870 1450
rect 980 1110 1040 1450
<< ndiff >>
rect 560 380 660 390
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 470 380
rect 530 370 700 380
rect 530 230 592 370
rect 638 230 700 370
rect 530 210 700 230
rect 760 210 810 380
rect 870 318 980 380
rect 870 272 902 318
rect 948 272 980 318
rect 870 210 980 272
rect 1040 318 1140 380
rect 1040 272 1072 318
rect 1118 272 1140 318
rect 1040 210 1140 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1110 470 1450
rect 530 1397 700 1450
rect 530 1163 592 1397
rect 638 1163 700 1397
rect 530 1110 700 1163
rect 760 1110 810 1450
rect 870 1397 980 1450
rect 870 1163 902 1397
rect 948 1163 980 1397
rect 870 1110 980 1163
rect 1040 1397 1140 1450
rect 1040 1163 1072 1397
rect 1118 1163 1140 1397
rect 1040 1110 1140 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 592 230 638 370
rect 902 272 948 318
rect 1072 272 1118 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 592 1163 638 1397
rect 902 1163 948 1397
rect 1072 1163 1118 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1020 1588 1170 1610
rect 1020 1542 1072 1588
rect 1118 1542 1170 1588
rect 1020 1520 1170 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1072 1542 1118 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 470 1450 530 1500
rect 700 1450 760 1500
rect 810 1450 870 1500
rect 980 1450 1040 1500
rect 190 540 250 1110
rect 360 800 420 1110
rect 310 773 420 800
rect 310 727 337 773
rect 383 727 420 773
rect 310 700 420 727
rect 470 930 530 1110
rect 470 903 610 930
rect 470 857 537 903
rect 583 857 610 903
rect 470 830 610 857
rect 190 513 350 540
rect 190 467 277 513
rect 323 490 350 513
rect 323 467 420 490
rect 190 430 420 467
rect 190 380 250 430
rect 360 380 420 430
rect 470 380 530 830
rect 700 800 760 1110
rect 810 1060 870 1110
rect 980 1060 1040 1110
rect 810 1000 1040 1060
rect 690 773 810 800
rect 690 727 737 773
rect 783 727 810 773
rect 690 700 810 727
rect 980 540 1040 1000
rect 580 520 680 540
rect 580 513 760 520
rect 580 467 607 513
rect 653 467 760 513
rect 870 513 1040 540
rect 870 490 897 513
rect 580 440 760 467
rect 700 380 760 440
rect 810 467 897 490
rect 943 467 1040 513
rect 810 440 1040 467
rect 810 380 870 440
rect 980 380 1040 440
rect 190 160 250 210
rect 360 160 420 210
rect 470 160 530 210
rect 700 160 760 210
rect 810 160 870 210
rect 980 160 1040 210
<< polycontact >>
rect 337 727 383 773
rect 537 857 583 903
rect 277 467 323 513
rect 737 727 783 773
rect 607 467 653 513
rect 897 467 943 513
<< metal1 >>
rect 0 1588 1240 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1072 1588
rect 1118 1542 1240 1588
rect 0 1520 1240 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 780 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 590 1397 640 1450
rect 590 1190 592 1397
rect 280 1110 330 1163
rect 580 1166 592 1190
rect 580 1114 584 1166
rect 638 1163 640 1397
rect 636 1114 640 1163
rect 580 1080 640 1114
rect 900 1397 950 1520
rect 900 1163 902 1397
rect 948 1163 950 1397
rect 900 1110 950 1163
rect 1070 1397 1120 1450
rect 1070 1163 1072 1397
rect 1118 1163 1120 1397
rect 1070 910 1120 1163
rect 510 903 1120 910
rect 510 857 537 903
rect 583 857 1120 903
rect 510 850 1120 857
rect 110 773 660 780
rect 110 727 337 773
rect 383 727 660 773
rect 110 720 660 727
rect 710 776 810 780
rect 710 724 734 776
rect 786 724 810 776
rect 710 720 810 724
rect 110 318 160 720
rect 600 520 660 720
rect 250 516 350 520
rect 250 464 274 516
rect 326 464 350 516
rect 250 460 350 464
rect 580 513 680 520
rect 580 467 607 513
rect 653 467 680 513
rect 580 460 680 467
rect 870 516 970 520
rect 870 464 894 516
rect 946 464 970 516
rect 870 460 970 464
rect 580 386 640 410
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 580 334 584 386
rect 636 370 640 386
rect 580 300 592 334
rect 280 140 330 272
rect 590 230 592 300
rect 638 230 640 370
rect 590 210 640 230
rect 900 318 950 380
rect 900 272 902 318
rect 948 272 950 318
rect 900 140 950 272
rect 1070 318 1120 850
rect 1070 272 1072 318
rect 1118 272 1120 318
rect 1070 210 1120 272
rect 0 118 1240 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1240 118
rect 0 0 1240 72
<< via1 >>
rect 584 1163 592 1166
rect 592 1163 636 1166
rect 584 1114 636 1163
rect 734 773 786 776
rect 734 727 737 773
rect 737 727 783 773
rect 783 727 786 773
rect 734 724 786 727
rect 274 513 326 516
rect 274 467 277 513
rect 277 467 323 513
rect 323 467 326 513
rect 274 464 326 467
rect 894 513 946 516
rect 894 467 897 513
rect 897 467 943 513
rect 943 467 946 513
rect 894 464 946 467
rect 584 370 636 386
rect 584 334 592 370
rect 592 334 636 370
<< metal2 >>
rect 580 1180 640 1210
rect 570 1166 650 1180
rect 570 1114 584 1166
rect 636 1114 650 1166
rect 570 1100 650 1114
rect 270 530 330 540
rect 260 516 340 530
rect 260 464 274 516
rect 326 464 340 516
rect 260 450 340 464
rect 270 260 330 450
rect 580 400 640 1100
rect 730 790 790 800
rect 720 776 800 790
rect 720 724 734 776
rect 786 724 800 776
rect 720 710 800 724
rect 560 386 660 400
rect 560 334 584 386
rect 636 334 660 386
rect 560 320 660 334
rect 730 260 790 710
rect 890 530 950 540
rect 880 520 960 530
rect 870 516 970 520
rect 870 464 894 516
rect 946 464 970 516
rect 870 460 970 464
rect 880 450 960 460
rect 890 440 950 450
rect 270 200 790 260
<< labels >>
rlabel via1 s 734 724 786 776 4 A
port 1 nsew signal input
rlabel via1 s 894 464 946 516 4 B
port 2 nsew signal input
rlabel via1 s 584 334 636 386 4 Y
port 3 nsew signal output
rlabel metal1 s 280 1110 330 1660 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 900 1110 950 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1520 1240 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 900 0 950 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1240 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 274 464 326 516 1 A
port 1 nsew signal input
rlabel metal2 s 270 200 330 540 1 A
port 1 nsew signal input
rlabel metal2 s 260 450 340 530 1 A
port 1 nsew signal input
rlabel metal2 s 270 200 790 260 1 A
port 1 nsew signal input
rlabel metal2 s 730 200 790 800 1 A
port 1 nsew signal input
rlabel metal2 s 720 710 800 790 1 A
port 1 nsew signal input
rlabel metal1 s 250 460 350 520 1 A
port 1 nsew signal input
rlabel metal1 s 710 720 810 780 1 A
port 1 nsew signal input
rlabel metal2 s 890 440 950 540 1 B
port 2 nsew signal input
rlabel metal2 s 880 450 960 530 1 B
port 2 nsew signal input
rlabel metal2 s 870 460 970 520 1 B
port 2 nsew signal input
rlabel metal1 s 870 460 970 520 1 B
port 2 nsew signal input
rlabel via1 s 584 1114 636 1166 1 Y
port 3 nsew signal output
rlabel metal2 s 580 320 640 1210 1 Y
port 3 nsew signal output
rlabel metal2 s 570 1100 650 1180 1 Y
port 3 nsew signal output
rlabel metal2 s 560 320 660 400 1 Y
port 3 nsew signal output
rlabel metal1 s 580 1080 640 1190 1 Y
port 3 nsew signal output
rlabel metal1 s 590 1080 640 1450 1 Y
port 3 nsew signal output
rlabel metal1 s 590 210 640 410 1 Y
port 3 nsew signal output
rlabel metal1 s 580 300 640 410 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1240 1660
string GDS_END 524418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 515772
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
