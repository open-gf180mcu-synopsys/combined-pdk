magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 440 1270
<< nmos >>
rect 190 210 250 380
<< pmos >>
rect 190 720 250 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 298 350 380
rect 250 252 282 298
rect 328 252 350 298
rect 250 210 350 252
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 350 1060
rect 250 773 282 1007
rect 328 773 350 1007
rect 250 720 350 773
<< ndiffc >>
rect 112 272 158 318
rect 282 252 328 298
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
<< psubdiffcont >>
rect 112 72 158 118
<< nsubdiffcont >>
rect 112 1152 158 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 190 670 250 720
rect 190 648 330 670
rect 190 602 262 648
rect 308 602 330 648
rect 190 580 330 602
rect 190 380 250 580
rect 190 160 250 210
<< polycontact >>
rect 262 602 308 648
<< metal1 >>
rect 0 1198 440 1270
rect 0 1152 112 1198
rect 158 1152 440 1198
rect 0 1130 440 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 650 330 773
rect 230 648 330 650
rect 230 602 262 648
rect 308 602 330 648
rect 230 600 330 602
rect 280 390 330 400
rect 260 386 360 390
rect 110 318 160 380
rect 260 334 284 386
rect 336 334 360 386
rect 260 330 360 334
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 298 330 330
rect 280 252 282 298
rect 328 252 330 298
rect 280 210 330 252
rect 0 118 440 140
rect 0 72 112 118
rect 158 72 440 118
rect 0 0 440 72
<< via1 >>
rect 284 334 336 386
<< metal2 >>
rect 260 386 360 400
rect 260 334 284 386
rect 336 334 360 386
rect 260 320 360 334
<< labels >>
rlabel via1 s 284 334 336 386 4 Y
port 1 nsew signal output
rlabel metal1 s 110 720 160 1270 4 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 1130 440 1270 1 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 0 440 140 1 VSS
port 3 nsew ground bidirectional abutment
rlabel metal2 s 260 320 360 400 1 Y
port 1 nsew signal output
rlabel metal1 s 280 210 330 400 1 Y
port 1 nsew signal output
rlabel metal1 s 260 330 360 390 1 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 440 1270
string GDS_END 372648
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 370094
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
