magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 460 1660
rect 580 1020 1560 1660
<< nmos >>
rect 200 210 260 380
rect 780 210 840 380
rect 960 210 1020 380
rect 1300 210 1360 380
<< pmos >>
rect 200 1110 260 1450
rect 780 1110 840 1450
rect 960 1110 1020 1450
rect 1300 1110 1360 1450
<< ndiff >>
rect 90 318 200 380
rect 90 272 117 318
rect 163 272 200 318
rect 90 210 200 272
rect 260 318 370 380
rect 260 272 297 318
rect 343 272 370 318
rect 260 210 370 272
rect 670 318 780 380
rect 670 272 697 318
rect 743 272 780 318
rect 670 210 780 272
rect 840 318 960 380
rect 840 272 877 318
rect 923 272 960 318
rect 840 210 960 272
rect 1020 318 1130 380
rect 1020 272 1057 318
rect 1103 272 1130 318
rect 1020 210 1130 272
rect 1190 318 1300 380
rect 1190 272 1217 318
rect 1263 272 1300 318
rect 1190 210 1300 272
rect 1360 318 1470 380
rect 1360 272 1397 318
rect 1443 272 1470 318
rect 1360 210 1470 272
<< pdiff >>
rect 90 1397 200 1450
rect 90 1163 117 1397
rect 163 1163 200 1397
rect 90 1110 200 1163
rect 260 1397 370 1450
rect 260 1163 297 1397
rect 343 1163 370 1397
rect 260 1110 370 1163
rect 670 1397 780 1450
rect 670 1163 697 1397
rect 743 1163 780 1397
rect 670 1110 780 1163
rect 840 1397 960 1450
rect 840 1163 877 1397
rect 923 1163 960 1397
rect 840 1110 960 1163
rect 1020 1397 1130 1450
rect 1020 1163 1057 1397
rect 1103 1163 1130 1397
rect 1020 1110 1130 1163
rect 1190 1397 1300 1450
rect 1190 1163 1217 1397
rect 1263 1163 1300 1397
rect 1190 1110 1300 1163
rect 1360 1397 1470 1450
rect 1360 1163 1397 1397
rect 1443 1163 1470 1397
rect 1360 1110 1470 1163
<< ndiffc >>
rect 117 272 163 318
rect 297 272 343 318
rect 697 272 743 318
rect 877 272 923 318
rect 1057 272 1103 318
rect 1217 272 1263 318
rect 1397 272 1443 318
<< pdiffc >>
rect 117 1163 163 1397
rect 297 1163 343 1397
rect 697 1163 743 1397
rect 877 1163 923 1397
rect 1057 1163 1103 1397
rect 1217 1163 1263 1397
rect 1397 1163 1443 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
rect 980 118 1130 140
rect 980 72 1032 118
rect 1078 72 1130 118
rect 980 50 1130 72
rect 1210 118 1360 140
rect 1210 72 1262 118
rect 1308 72 1360 118
rect 1210 50 1360 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 640 1588 790 1610
rect 640 1542 692 1588
rect 738 1542 790 1588
rect 640 1520 790 1542
rect 870 1588 1020 1610
rect 870 1542 922 1588
rect 968 1542 1020 1588
rect 870 1520 1020 1542
rect 1100 1588 1250 1610
rect 1100 1542 1152 1588
rect 1198 1542 1250 1588
rect 1100 1520 1250 1542
rect 1330 1588 1480 1610
rect 1330 1542 1382 1588
rect 1428 1542 1480 1588
rect 1330 1520 1480 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
rect 1032 72 1078 118
rect 1262 72 1308 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 692 1542 738 1588
rect 922 1542 968 1588
rect 1152 1542 1198 1588
rect 1382 1542 1428 1588
<< polysilicon >>
rect 200 1450 260 1500
rect 780 1450 840 1500
rect 960 1450 1020 1500
rect 1300 1450 1360 1500
rect 200 540 260 1110
rect 780 900 840 1110
rect 960 1060 1020 1110
rect 1300 1060 1360 1110
rect 910 1038 1020 1060
rect 910 992 932 1038
rect 978 992 1020 1038
rect 910 980 1020 992
rect 1230 1038 1360 1060
rect 1230 992 1252 1038
rect 1298 992 1360 1038
rect 910 970 1000 980
rect 1230 970 1360 992
rect 960 900 1050 910
rect 780 888 1050 900
rect 780 842 982 888
rect 1028 842 1050 888
rect 780 840 1050 842
rect 960 820 1050 840
rect 900 658 1020 680
rect 900 612 932 658
rect 978 612 1020 658
rect 900 590 1020 612
rect 120 518 260 540
rect 120 472 152 518
rect 198 472 260 518
rect 120 450 260 472
rect 200 380 260 450
rect 780 518 900 540
rect 780 472 832 518
rect 878 472 900 518
rect 780 450 900 472
rect 780 380 840 450
rect 960 380 1020 590
rect 1300 380 1360 970
rect 200 160 260 210
rect 780 160 840 210
rect 960 160 1020 210
rect 1300 160 1360 210
<< polycontact >>
rect 932 992 978 1038
rect 1252 992 1298 1038
rect 982 842 1028 888
rect 932 612 978 658
rect 152 472 198 518
rect 832 472 878 518
<< metal1 >>
rect 0 1588 460 1660
rect 0 1542 112 1588
rect 158 1542 460 1588
rect 0 1520 460 1542
rect 580 1588 1560 1660
rect 580 1542 692 1588
rect 738 1542 922 1588
rect 968 1542 1152 1588
rect 1198 1542 1382 1588
rect 1428 1542 1560 1588
rect 580 1520 1560 1542
rect 110 1397 170 1520
rect 110 1163 117 1397
rect 163 1163 170 1397
rect 110 1110 170 1163
rect 290 1397 350 1450
rect 290 1163 297 1397
rect 343 1163 350 1397
rect 290 660 350 1163
rect 690 1397 750 1450
rect 690 1163 697 1397
rect 743 1163 750 1397
rect 690 1040 750 1163
rect 870 1397 930 1520
rect 870 1163 877 1397
rect 923 1163 930 1397
rect 870 1110 930 1163
rect 1050 1397 1110 1450
rect 1050 1163 1057 1397
rect 1103 1163 1110 1397
rect 910 1040 1000 1060
rect 690 1038 1000 1040
rect 690 1036 932 1038
rect 690 984 924 1036
rect 978 992 1000 1038
rect 976 984 1000 992
rect 690 980 1000 984
rect 270 656 370 660
rect 270 604 294 656
rect 346 604 370 656
rect 270 600 370 604
rect 120 518 220 520
rect 120 516 152 518
rect 120 464 144 516
rect 198 472 220 518
rect 196 464 220 472
rect 120 460 220 464
rect 110 318 170 380
rect 110 272 117 318
rect 163 272 170 318
rect 110 140 170 272
rect 290 318 350 600
rect 290 272 297 318
rect 343 272 350 318
rect 290 210 350 272
rect 690 318 750 980
rect 910 970 1000 980
rect 1050 910 1110 1163
rect 1210 1397 1270 1520
rect 1210 1163 1217 1397
rect 1263 1163 1270 1397
rect 1210 1110 1270 1163
rect 1390 1397 1450 1450
rect 1390 1163 1397 1397
rect 1443 1163 1450 1397
rect 1220 1038 1320 1040
rect 1220 1036 1252 1038
rect 1220 984 1244 1036
rect 1298 992 1320 1038
rect 1296 984 1320 992
rect 1220 980 1320 984
rect 1390 910 1450 1163
rect 960 888 1110 910
rect 960 842 982 888
rect 1028 842 1110 888
rect 1380 906 1460 910
rect 1380 854 1394 906
rect 1446 854 1460 906
rect 1380 850 1460 854
rect 960 820 1110 842
rect 900 658 1000 660
rect 900 656 932 658
rect 900 604 924 656
rect 978 612 1000 658
rect 976 604 1000 612
rect 900 600 1000 604
rect 800 518 900 520
rect 800 516 832 518
rect 800 464 824 516
rect 878 472 900 518
rect 876 464 900 472
rect 800 460 900 464
rect 690 272 697 318
rect 743 272 750 318
rect 690 210 750 272
rect 870 318 930 380
rect 870 272 877 318
rect 923 272 930 318
rect 870 140 930 272
rect 1050 318 1110 820
rect 1050 272 1057 318
rect 1103 272 1110 318
rect 1050 210 1110 272
rect 1210 318 1270 380
rect 1210 272 1217 318
rect 1263 272 1270 318
rect 1210 140 1270 272
rect 1390 318 1450 850
rect 1390 272 1397 318
rect 1443 272 1450 318
rect 1390 210 1450 272
rect 0 118 1560 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1032 118
rect 1078 72 1262 118
rect 1308 72 1560 118
rect 0 0 1560 72
<< via1 >>
rect 924 992 932 1036
rect 932 992 976 1036
rect 924 984 976 992
rect 294 604 346 656
rect 144 472 152 516
rect 152 472 196 516
rect 144 464 196 472
rect 1244 992 1252 1036
rect 1252 992 1296 1036
rect 1244 984 1296 992
rect 1394 854 1446 906
rect 924 612 932 656
rect 932 612 976 656
rect 924 604 976 612
rect 824 472 832 516
rect 832 472 876 516
rect 824 464 876 472
<< metal2 >>
rect 910 1040 990 1050
rect 1220 1040 1320 1050
rect 900 1036 1320 1040
rect 900 984 924 1036
rect 976 984 1244 1036
rect 1296 984 1320 1036
rect 900 980 1320 984
rect 910 970 990 980
rect 1220 970 1320 980
rect 1370 906 1470 920
rect 1370 854 1394 906
rect 1446 854 1470 906
rect 1370 840 1470 854
rect 270 660 370 670
rect 900 660 1000 670
rect 270 656 1000 660
rect 270 604 294 656
rect 346 604 924 656
rect 976 604 1000 656
rect 270 600 1000 604
rect 270 590 370 600
rect 900 590 1000 600
rect 120 520 220 530
rect 800 520 900 530
rect 120 516 900 520
rect 120 464 144 516
rect 196 464 824 516
rect 876 464 900 516
rect 120 460 900 464
rect 120 450 220 460
rect 800 450 900 460
<< labels >>
rlabel via1 s 824 464 876 516 4 A
port 1 nsew signal input
rlabel via1 s 1394 854 1446 906 4 Y
port 2 nsew signal output
rlabel metal1 s 870 1110 930 1660 4 VDDH
port 3 nsew power bidirectional
rlabel metal1 s 110 1110 170 1660 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 110 0 170 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 1520 460 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1210 1110 1270 1660 1 VDDH
port 3 nsew power bidirectional
rlabel metal1 s 580 1520 1560 1660 1 VDDH
port 3 nsew power bidirectional
rlabel metal1 s 870 0 930 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1210 0 1270 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1560 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 144 464 196 516 1 A
port 1 nsew signal input
rlabel metal2 s 120 450 220 530 1 A
port 1 nsew signal input
rlabel metal2 s 120 460 900 520 1 A
port 1 nsew signal input
rlabel metal2 s 800 450 900 530 1 A
port 1 nsew signal input
rlabel metal1 s 120 460 220 520 1 A
port 1 nsew signal input
rlabel metal1 s 800 460 900 520 1 A
port 1 nsew signal input
rlabel metal2 s 1370 840 1470 920 1 Y
port 2 nsew signal output
rlabel metal1 s 1390 210 1450 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 1380 850 1460 910 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1560 1660
string GDS_END 457638
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 447838
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
