magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 2600 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 520 210 580 380
rect 690 210 750 380
rect 800 210 860 380
rect 970 210 1030 380
rect 1080 210 1140 380
rect 1250 210 1310 380
rect 1360 210 1420 380
rect 1530 210 1590 380
rect 1850 210 1910 380
rect 2170 210 2230 380
rect 2340 210 2400 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 520 1110 580 1450
rect 690 1110 750 1450
rect 800 1110 860 1450
rect 970 1110 1030 1450
rect 1080 1110 1140 1450
rect 1250 1110 1310 1450
rect 1360 1110 1420 1450
rect 1530 1110 1590 1450
rect 1850 1110 1910 1450
rect 2170 1110 2230 1450
rect 2340 1110 2400 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 520 380
rect 580 318 690 380
rect 580 272 612 318
rect 658 272 690 318
rect 580 210 690 272
rect 750 210 800 380
rect 860 278 970 380
rect 860 232 892 278
rect 938 232 970 278
rect 860 210 970 232
rect 1030 210 1080 380
rect 1140 318 1250 380
rect 1140 272 1172 318
rect 1218 272 1250 318
rect 1140 210 1250 272
rect 1310 210 1360 380
rect 1420 318 1530 380
rect 1420 272 1452 318
rect 1498 272 1530 318
rect 1420 210 1530 272
rect 1590 318 1690 380
rect 1590 272 1622 318
rect 1668 272 1690 318
rect 1590 210 1690 272
rect 1750 283 1850 380
rect 1750 237 1772 283
rect 1818 237 1850 283
rect 1750 210 1850 237
rect 1910 318 2010 380
rect 1910 272 1942 318
rect 1988 272 2010 318
rect 1910 210 2010 272
rect 2070 318 2170 380
rect 2070 272 2092 318
rect 2138 272 2170 318
rect 2070 210 2170 272
rect 2230 318 2340 380
rect 2230 272 2262 318
rect 2308 272 2340 318
rect 2230 210 2340 272
rect 2400 318 2500 380
rect 2400 272 2432 318
rect 2478 272 2500 318
rect 2400 210 2500 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1110 520 1450
rect 580 1397 690 1450
rect 580 1163 612 1397
rect 658 1163 690 1397
rect 580 1110 690 1163
rect 750 1110 800 1450
rect 860 1397 970 1450
rect 860 1163 892 1397
rect 938 1163 970 1397
rect 860 1110 970 1163
rect 1030 1110 1080 1450
rect 1140 1425 1250 1450
rect 1140 1285 1172 1425
rect 1218 1285 1250 1425
rect 1140 1110 1250 1285
rect 1310 1110 1360 1450
rect 1420 1425 1530 1450
rect 1420 1285 1452 1425
rect 1498 1285 1530 1425
rect 1420 1110 1530 1285
rect 1590 1397 1690 1450
rect 1590 1163 1622 1397
rect 1668 1163 1690 1397
rect 1590 1110 1690 1163
rect 1750 1397 1850 1450
rect 1750 1163 1772 1397
rect 1818 1163 1850 1397
rect 1750 1110 1850 1163
rect 1910 1397 2010 1450
rect 1910 1163 1942 1397
rect 1988 1163 2010 1397
rect 1910 1110 2010 1163
rect 2070 1397 2170 1450
rect 2070 1163 2092 1397
rect 2138 1163 2170 1397
rect 2070 1110 2170 1163
rect 2230 1397 2340 1450
rect 2230 1163 2262 1397
rect 2308 1163 2340 1397
rect 2230 1110 2340 1163
rect 2400 1397 2500 1450
rect 2400 1163 2432 1397
rect 2478 1163 2500 1397
rect 2400 1110 2500 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 612 272 658 318
rect 892 232 938 278
rect 1172 272 1218 318
rect 1452 272 1498 318
rect 1622 272 1668 318
rect 1772 237 1818 283
rect 1942 272 1988 318
rect 2092 272 2138 318
rect 2262 272 2308 318
rect 2432 272 2478 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 612 1163 658 1397
rect 892 1163 938 1397
rect 1172 1285 1218 1425
rect 1452 1285 1498 1425
rect 1622 1163 1668 1397
rect 1772 1163 1818 1397
rect 1942 1163 1988 1397
rect 2092 1163 2138 1397
rect 2262 1163 2308 1397
rect 2432 1163 2478 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1020 1588 1170 1610
rect 1020 1542 1072 1588
rect 1118 1542 1170 1588
rect 1020 1520 1170 1542
rect 1260 1588 1410 1610
rect 1260 1542 1312 1588
rect 1358 1542 1410 1588
rect 1260 1520 1410 1542
rect 1500 1588 1650 1610
rect 1500 1542 1552 1588
rect 1598 1542 1650 1588
rect 1500 1520 1650 1542
rect 1740 1588 1890 1610
rect 1740 1542 1792 1588
rect 1838 1542 1890 1588
rect 1740 1520 1890 1542
rect 1980 1588 2130 1610
rect 1980 1542 2032 1588
rect 2078 1542 2130 1588
rect 1980 1520 2130 1542
rect 2220 1588 2370 1610
rect 2220 1542 2272 1588
rect 2318 1542 2370 1588
rect 2220 1520 2370 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1072 1542 1118 1588
rect 1312 1542 1358 1588
rect 1552 1542 1598 1588
rect 1792 1542 1838 1588
rect 2032 1542 2078 1588
rect 2272 1542 2318 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 520 1450 580 1500
rect 690 1450 750 1500
rect 800 1450 860 1500
rect 970 1450 1030 1500
rect 1080 1450 1140 1500
rect 1250 1450 1310 1500
rect 1360 1450 1420 1500
rect 1530 1450 1590 1500
rect 1850 1450 1910 1500
rect 2170 1450 2230 1500
rect 2340 1450 2400 1500
rect 190 930 250 1110
rect 190 903 310 930
rect 190 857 237 903
rect 283 857 310 903
rect 190 830 310 857
rect 190 380 250 830
rect 360 800 420 1110
rect 520 930 580 1110
rect 520 903 620 930
rect 520 857 547 903
rect 593 857 620 903
rect 520 830 620 857
rect 360 773 480 800
rect 360 727 407 773
rect 453 727 480 773
rect 360 700 480 727
rect 360 380 420 700
rect 690 660 750 1110
rect 800 1060 860 1110
rect 970 1060 1030 1110
rect 800 1033 1030 1060
rect 800 990 837 1033
rect 810 987 837 990
rect 883 990 1030 1033
rect 883 987 910 990
rect 810 940 910 987
rect 1080 660 1140 1110
rect 1250 930 1310 1110
rect 1210 903 1310 930
rect 1210 857 1237 903
rect 1283 857 1310 903
rect 1210 830 1310 857
rect 1360 800 1420 1110
rect 1530 930 1590 1110
rect 1530 903 1630 930
rect 1530 857 1557 903
rect 1603 857 1630 903
rect 1530 830 1630 857
rect 1350 773 1460 800
rect 1350 727 1377 773
rect 1423 727 1460 773
rect 1350 700 1460 727
rect 1210 660 1310 670
rect 520 643 1310 660
rect 520 600 1237 643
rect 520 380 580 600
rect 1210 597 1237 600
rect 1283 597 1310 643
rect 1210 570 1310 597
rect 650 513 750 540
rect 810 520 910 540
rect 650 467 677 513
rect 723 467 750 513
rect 650 440 750 467
rect 690 380 750 440
rect 800 513 1030 520
rect 800 467 837 513
rect 883 467 1030 513
rect 800 440 1030 467
rect 800 380 860 440
rect 970 380 1030 440
rect 1080 503 1180 530
rect 1080 457 1107 503
rect 1153 457 1180 503
rect 1080 430 1180 457
rect 1080 380 1140 430
rect 1250 380 1310 570
rect 1360 380 1420 700
rect 1530 380 1590 830
rect 1850 670 1910 1110
rect 2170 670 2230 1110
rect 2340 930 2400 1110
rect 2280 903 2400 930
rect 2280 857 2307 903
rect 2353 857 2400 903
rect 2280 830 2400 857
rect 1790 643 1910 670
rect 1790 597 1817 643
rect 1863 597 1910 643
rect 1790 570 1910 597
rect 2110 643 2230 670
rect 2110 597 2157 643
rect 2203 597 2230 643
rect 2110 570 2230 597
rect 1850 380 1910 570
rect 2170 380 2230 570
rect 2340 380 2400 830
rect 190 160 250 210
rect 360 160 420 210
rect 520 160 580 210
rect 690 160 750 210
rect 800 160 860 210
rect 970 160 1030 210
rect 1080 160 1140 210
rect 1250 160 1310 210
rect 1360 160 1420 210
rect 1530 160 1590 210
rect 1850 160 1910 210
rect 2170 160 2230 210
rect 2340 160 2400 210
<< polycontact >>
rect 237 857 283 903
rect 547 857 593 903
rect 407 727 453 773
rect 837 987 883 1033
rect 1237 857 1283 903
rect 1557 857 1603 903
rect 1377 727 1423 773
rect 1237 597 1283 643
rect 677 467 723 513
rect 837 467 883 513
rect 1107 457 1153 503
rect 2307 857 2353 903
rect 1817 597 1863 643
rect 2157 597 2203 643
<< metal1 >>
rect 0 1588 2600 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1072 1588
rect 1118 1542 1312 1588
rect 1358 1542 1552 1588
rect 1598 1542 1792 1588
rect 1838 1542 2032 1588
rect 2078 1542 2272 1588
rect 2318 1542 2600 1588
rect 0 1520 2600 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 540 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 610 1397 660 1450
rect 610 1163 612 1397
rect 658 1163 660 1397
rect 610 1060 660 1163
rect 890 1397 940 1520
rect 890 1163 892 1397
rect 938 1163 940 1397
rect 1170 1425 1220 1450
rect 1170 1285 1172 1425
rect 1218 1285 1220 1425
rect 1170 1260 1220 1285
rect 1450 1425 1500 1520
rect 1450 1285 1452 1425
rect 1498 1285 1500 1425
rect 1450 1260 1500 1285
rect 1620 1397 1670 1450
rect 890 1110 940 1163
rect 990 1210 1220 1260
rect 280 1010 660 1060
rect 810 1033 910 1040
rect 280 910 330 1010
rect 810 987 837 1033
rect 883 987 910 1033
rect 810 980 910 987
rect 210 903 330 910
rect 210 857 237 903
rect 283 857 330 903
rect 210 850 330 857
rect 520 906 750 910
rect 520 903 674 906
rect 520 857 547 903
rect 593 857 674 903
rect 520 854 674 857
rect 726 854 750 906
rect 520 850 750 854
rect 100 516 160 540
rect 100 464 104 516
rect 156 464 160 516
rect 280 520 330 850
rect 380 776 480 780
rect 380 724 404 776
rect 456 724 480 776
rect 380 720 480 724
rect 670 520 730 850
rect 830 520 890 980
rect 990 760 1040 1210
rect 1620 1163 1622 1397
rect 1668 1163 1670 1397
rect 1340 1036 1440 1040
rect 1340 984 1364 1036
rect 1416 984 1440 1036
rect 1340 980 1440 984
rect 1620 1020 1670 1163
rect 1770 1397 1820 1520
rect 1770 1163 1772 1397
rect 1818 1163 1820 1397
rect 1770 1110 1820 1163
rect 1940 1397 1990 1450
rect 1940 1163 1942 1397
rect 1988 1163 1990 1397
rect 980 710 1040 760
rect 1100 906 1310 910
rect 1100 854 1234 906
rect 1286 854 1310 906
rect 1100 850 1310 854
rect 280 470 480 520
rect 100 440 160 464
rect 110 318 160 440
rect 400 380 480 470
rect 650 513 750 520
rect 650 467 677 513
rect 723 467 750 513
rect 650 460 750 467
rect 810 516 910 520
rect 810 464 834 516
rect 886 464 910 516
rect 810 460 910 464
rect 980 390 1030 710
rect 1100 510 1160 850
rect 1360 780 1420 980
rect 1620 970 1780 1020
rect 1530 906 1630 910
rect 1530 854 1554 906
rect 1606 854 1630 906
rect 1530 850 1630 854
rect 1720 780 1780 970
rect 1350 776 1460 780
rect 1350 724 1374 776
rect 1426 724 1460 776
rect 1350 720 1460 724
rect 1620 730 1780 780
rect 1360 710 1440 720
rect 1210 646 1310 650
rect 1210 594 1234 646
rect 1286 594 1310 646
rect 1210 590 1310 594
rect 1620 646 1680 730
rect 1810 650 1870 670
rect 1940 650 1990 1163
rect 2090 1397 2140 1450
rect 2090 1163 2092 1397
rect 2138 1163 2140 1397
rect 2090 910 2140 1163
rect 2260 1397 2310 1520
rect 2260 1163 2262 1397
rect 2308 1163 2310 1397
rect 2260 1110 2310 1163
rect 2430 1397 2480 1450
rect 2430 1163 2432 1397
rect 2478 1163 2480 1397
rect 2430 1050 2480 1163
rect 2430 1036 2530 1050
rect 2430 984 2454 1036
rect 2506 984 2530 1036
rect 2430 980 2530 984
rect 2430 970 2520 980
rect 2090 906 2380 910
rect 2090 854 2304 906
rect 2356 854 2380 906
rect 2090 850 2380 854
rect 1620 594 1624 646
rect 1676 594 1680 646
rect 1620 570 1680 594
rect 1790 643 1890 650
rect 1790 597 1817 643
rect 1863 597 1890 643
rect 1790 590 1890 597
rect 1940 646 2230 650
rect 1940 594 2154 646
rect 2206 594 2230 646
rect 1940 590 2230 594
rect 1080 503 1180 510
rect 1080 457 1107 503
rect 1153 457 1180 503
rect 1080 450 1180 457
rect 980 386 1250 390
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 400 330 660 380
rect 980 340 1174 386
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 610 318 660 330
rect 610 272 612 318
rect 658 272 660 318
rect 1170 334 1174 340
rect 1226 334 1250 386
rect 1170 330 1250 334
rect 1170 318 1220 330
rect 610 210 660 272
rect 890 278 940 300
rect 890 232 892 278
rect 938 232 940 278
rect 890 140 940 232
rect 1170 272 1172 318
rect 1218 272 1220 318
rect 1170 210 1220 272
rect 1450 318 1500 380
rect 1450 272 1452 318
rect 1498 272 1500 318
rect 1450 140 1500 272
rect 1620 318 1670 570
rect 1810 420 1870 590
rect 1790 416 1890 420
rect 1790 364 1814 416
rect 1866 364 1890 416
rect 1790 360 1890 364
rect 1620 272 1622 318
rect 1668 272 1670 318
rect 1940 318 1990 590
rect 2310 480 2360 850
rect 1620 210 1670 272
rect 1770 283 1820 310
rect 1770 237 1772 283
rect 1818 237 1820 283
rect 1770 140 1820 237
rect 1940 272 1942 318
rect 1988 272 1990 318
rect 1940 210 1990 272
rect 2090 430 2360 480
rect 2090 318 2140 430
rect 2090 272 2092 318
rect 2138 272 2140 318
rect 2090 210 2140 272
rect 2260 318 2310 380
rect 2260 272 2262 318
rect 2308 272 2310 318
rect 2260 140 2310 272
rect 2430 318 2480 970
rect 2430 272 2432 318
rect 2478 272 2480 318
rect 2430 210 2480 272
rect 0 118 2600 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2600 118
rect 0 0 2600 72
<< via1 >>
rect 674 854 726 906
rect 104 464 156 516
rect 404 773 456 776
rect 404 727 407 773
rect 407 727 453 773
rect 453 727 456 773
rect 404 724 456 727
rect 1364 984 1416 1036
rect 1234 903 1286 906
rect 1234 857 1237 903
rect 1237 857 1283 903
rect 1283 857 1286 903
rect 1234 854 1286 857
rect 834 513 886 516
rect 834 467 837 513
rect 837 467 883 513
rect 883 467 886 513
rect 834 464 886 467
rect 1554 903 1606 906
rect 1554 857 1557 903
rect 1557 857 1603 903
rect 1603 857 1606 903
rect 1554 854 1606 857
rect 1374 773 1426 776
rect 1374 727 1377 773
rect 1377 727 1423 773
rect 1423 727 1426 773
rect 1374 724 1426 727
rect 1234 643 1286 646
rect 1234 597 1237 643
rect 1237 597 1283 643
rect 1283 597 1286 643
rect 1234 594 1286 597
rect 2454 984 2506 1036
rect 2304 903 2356 906
rect 2304 857 2307 903
rect 2307 857 2353 903
rect 2353 857 2356 903
rect 2304 854 2356 857
rect 1624 594 1676 646
rect 2154 643 2206 646
rect 2154 597 2157 643
rect 2157 597 2203 643
rect 2203 597 2206 643
rect 2154 594 2206 597
rect 1174 334 1226 386
rect 1814 364 1866 416
<< metal2 >>
rect 1350 1040 1430 1050
rect 2440 1040 2520 1050
rect 1340 1036 1980 1040
rect 1340 984 1364 1036
rect 1416 984 1980 1036
rect 1340 980 1980 984
rect 2430 1036 2530 1040
rect 2430 984 2454 1036
rect 2506 984 2530 1036
rect 2430 980 2530 984
rect 1350 970 1430 980
rect 650 910 740 920
rect 1210 910 1310 920
rect 1540 910 1620 920
rect 650 906 1630 910
rect 650 854 674 906
rect 726 854 1234 906
rect 1286 854 1554 906
rect 1606 854 1630 906
rect 650 850 1630 854
rect 650 840 740 850
rect 1210 840 1310 850
rect 1540 840 1620 850
rect 380 780 480 790
rect 1360 780 1440 790
rect 350 776 510 780
rect 350 724 404 776
rect 456 724 510 776
rect 350 720 510 724
rect 1350 776 1450 780
rect 1350 724 1374 776
rect 1426 724 1450 776
rect 1350 720 1450 724
rect 380 710 480 720
rect 1360 710 1440 720
rect 1220 650 1300 660
rect 1610 650 1690 660
rect 1920 650 1980 980
rect 2440 970 2520 980
rect 2290 910 2370 920
rect 2280 906 2380 910
rect 2280 854 2304 906
rect 2356 854 2380 906
rect 2280 850 2380 854
rect 2290 840 2370 850
rect 2140 650 2220 660
rect 1210 646 1710 650
rect 1210 594 1234 646
rect 1286 594 1624 646
rect 1676 594 1710 646
rect 1210 590 1710 594
rect 1920 646 2230 650
rect 1920 594 2154 646
rect 2206 594 2230 646
rect 1920 590 2230 594
rect 1220 580 1300 590
rect 1610 580 1690 590
rect 2140 580 2220 590
rect 90 520 170 530
rect 820 520 900 530
rect 80 516 910 520
rect 80 464 104 516
rect 156 464 834 516
rect 886 464 910 516
rect 80 460 910 464
rect 90 450 170 460
rect 820 450 900 460
rect 1800 420 1880 430
rect 1700 416 1890 420
rect 1160 390 1240 400
rect 1700 390 1814 416
rect 1150 386 1814 390
rect 1150 334 1174 386
rect 1226 364 1814 386
rect 1866 364 1890 416
rect 1226 360 1890 364
rect 1226 350 1880 360
rect 1226 334 1760 350
rect 1150 330 1760 334
rect 1160 320 1240 330
<< labels >>
rlabel via1 s 404 724 456 776 4 D
port 1 nsew signal input
rlabel via1 s 2454 984 2506 1036 4 Q
port 2 nsew signal output
rlabel via1 s 2304 854 2356 906 4 QN
port 3 nsew signal output
rlabel via1 s 1554 854 1606 906 4 CLK
port 4 nsew clock input
rlabel metal1 s 280 1110 330 1660 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 890 1110 940 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1450 1260 1500 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1770 1110 1820 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2260 1110 2310 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1520 2600 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 890 0 940 300 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1450 0 1500 380 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1770 0 1820 310 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2260 0 2310 380 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2600 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel via1 s 1234 854 1286 906 1 CLK
port 4 nsew clock input
rlabel via1 s 674 854 726 906 1 CLK
port 4 nsew clock input
rlabel metal2 s 650 840 740 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 1210 840 1310 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 1540 840 1620 920 1 CLK
port 4 nsew clock input
rlabel metal2 s 650 850 1630 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 670 460 730 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 650 460 750 520 1 CLK
port 4 nsew clock input
rlabel metal1 s 520 850 750 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1100 450 1160 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1080 450 1180 510 1 CLK
port 4 nsew clock input
rlabel metal1 s 1100 850 1310 910 1 CLK
port 4 nsew clock input
rlabel metal1 s 1530 850 1630 910 1 CLK
port 4 nsew clock input
rlabel metal2 s 380 710 480 790 1 D
port 1 nsew signal input
rlabel metal2 s 350 720 510 780 1 D
port 1 nsew signal input
rlabel metal1 s 380 720 480 780 1 D
port 1 nsew signal input
rlabel metal2 s 2440 970 2520 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 2430 980 2530 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 210 2480 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 970 2520 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 980 2530 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 2290 840 2370 920 1 QN
port 3 nsew signal output
rlabel metal2 s 2280 850 2380 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 210 2140 480 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 850 2140 1450 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 430 2360 480 1 QN
port 3 nsew signal output
rlabel metal1 s 2310 430 2360 910 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 850 2380 910 1 QN
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2600 1660
string GDS_END 190270
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 170000
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
