magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 960 1660
<< nmos >>
rect 190 210 250 380
rect 530 210 590 380
rect 700 210 760 380
<< pmos >>
rect 190 1110 250 1450
rect 530 1110 590 1450
rect 700 1110 760 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 430 318 530 380
rect 430 272 452 318
rect 498 272 530 318
rect 430 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 318 860 380
rect 760 272 792 318
rect 838 272 860 318
rect 760 210 860 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 350 1450
rect 250 1163 282 1397
rect 328 1163 350 1397
rect 250 1110 350 1163
rect 430 1397 530 1450
rect 430 1163 452 1397
rect 498 1163 530 1397
rect 430 1110 530 1163
rect 590 1397 700 1450
rect 590 1163 622 1397
rect 668 1163 700 1397
rect 590 1110 700 1163
rect 760 1397 860 1450
rect 760 1163 792 1397
rect 838 1163 860 1397
rect 760 1110 860 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 792 272 838 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 452 1163 498 1397
rect 622 1163 668 1397
rect 792 1163 838 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 530 1450 590 1500
rect 700 1450 760 1500
rect 190 1080 250 1110
rect 530 1080 590 1110
rect 190 1030 590 1080
rect 190 670 250 1030
rect 300 910 400 940
rect 700 910 760 1110
rect 300 903 760 910
rect 300 857 327 903
rect 373 857 760 903
rect 300 850 760 857
rect 300 820 400 850
rect 120 650 250 670
rect 120 648 760 650
rect 120 602 142 648
rect 188 602 760 648
rect 120 600 760 602
rect 120 580 250 600
rect 190 380 250 580
rect 300 513 400 550
rect 300 467 327 513
rect 373 510 400 513
rect 373 467 590 510
rect 300 460 590 467
rect 300 430 400 460
rect 530 380 590 460
rect 700 380 760 600
rect 190 160 250 210
rect 530 160 590 210
rect 700 160 760 210
<< polycontact >>
rect 327 857 373 903
rect 142 602 188 648
rect 327 467 373 513
<< metal1 >>
rect 0 1588 960 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 960 1588
rect 0 1520 960 1542
rect 110 1397 160 1520
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1110 160 1163
rect 280 1397 330 1450
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 910 330 1163
rect 450 1397 500 1450
rect 450 1163 452 1397
rect 498 1163 500 1397
rect 280 903 400 910
rect 280 857 327 903
rect 373 857 400 903
rect 280 850 400 857
rect 110 648 210 650
rect 110 646 142 648
rect 110 594 134 646
rect 188 602 210 648
rect 186 594 210 602
rect 110 590 210 594
rect 280 520 330 850
rect 450 790 500 1163
rect 620 1397 670 1450
rect 620 1163 622 1397
rect 668 1163 670 1397
rect 620 1050 670 1163
rect 790 1397 840 1450
rect 790 1163 792 1397
rect 838 1163 840 1397
rect 600 1036 700 1050
rect 600 984 624 1036
rect 676 984 700 1036
rect 600 970 700 984
rect 450 776 570 790
rect 450 724 494 776
rect 546 724 570 776
rect 450 710 570 724
rect 280 513 400 520
rect 280 467 327 513
rect 373 467 400 513
rect 280 460 400 467
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 460
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 450 318 500 710
rect 450 272 452 318
rect 498 272 500 318
rect 450 210 500 272
rect 620 318 670 970
rect 790 920 840 1163
rect 750 906 850 920
rect 750 854 774 906
rect 826 854 850 906
rect 750 840 850 854
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 790 318 840 840
rect 790 272 792 318
rect 838 272 840 318
rect 790 210 840 272
rect 0 118 960 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 960 118
rect 0 0 960 72
<< via1 >>
rect 134 602 142 646
rect 142 602 186 646
rect 134 594 186 602
rect 624 984 676 1036
rect 494 724 546 776
rect 774 854 826 906
<< metal2 >>
rect 600 1036 700 1050
rect 600 984 624 1036
rect 676 984 700 1036
rect 600 970 700 984
rect 750 906 850 920
rect 750 854 774 906
rect 826 854 850 906
rect 750 840 850 854
rect 470 776 570 790
rect 470 724 494 776
rect 546 724 570 776
rect 470 710 570 724
rect 110 646 210 660
rect 110 594 134 646
rect 186 594 210 646
rect 110 580 210 594
<< labels >>
rlabel via1 s 494 724 546 776 4 A
port 1 nsew signal input
rlabel via1 s 774 854 826 906 4 B
port 2 nsew signal input
rlabel via1 s 624 984 676 1036 4 Y
port 3 nsew signal output
rlabel via1 s 134 594 186 646 4 Sel
port 4 nsew signal output
rlabel metal1 s 110 1110 160 1660 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 1520 960 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 0 960 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 470 710 570 790 1 A
port 1 nsew signal input
rlabel metal1 s 450 210 500 1450 1 A
port 1 nsew signal input
rlabel metal1 s 450 710 570 790 1 A
port 1 nsew signal input
rlabel metal2 s 750 840 850 920 1 B
port 2 nsew signal input
rlabel metal1 s 790 210 840 1450 1 B
port 2 nsew signal input
rlabel metal1 s 750 840 850 920 1 B
port 2 nsew signal input
rlabel metal2 s 110 580 210 660 1 Sel
port 4 nsew signal output
rlabel metal1 s 110 590 210 650 1 Sel
port 4 nsew signal output
rlabel metal2 s 600 970 700 1050 1 Y
port 3 nsew signal output
rlabel metal1 s 620 210 670 1450 1 Y
port 3 nsew signal output
rlabel metal1 s 600 970 700 1050 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 960 1660
string GDS_END 464340
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 457702
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
