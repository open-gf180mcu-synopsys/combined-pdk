magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 3160 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
rect 870 210 930 380
rect 1040 210 1100 380
rect 1210 210 1270 380
rect 1380 210 1440 380
rect 1550 210 1610 380
rect 1720 210 1780 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2400 210 2460 380
rect 2570 210 2630 380
rect 2740 210 2800 380
rect 2910 210 2970 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 530 1110 590 1450
rect 700 1110 760 1450
rect 870 1110 930 1450
rect 1040 1110 1100 1450
rect 1210 1110 1270 1450
rect 1380 1110 1440 1450
rect 1550 1110 1610 1450
rect 1720 1110 1780 1450
rect 1890 1110 1950 1450
rect 2060 1110 2120 1450
rect 2230 1110 2290 1450
rect 2400 1110 2460 1450
rect 2570 1110 2630 1450
rect 2740 1110 2800 1450
rect 2910 1110 2970 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 318 530 380
rect 420 272 452 318
rect 498 272 530 318
rect 420 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 318 870 380
rect 760 272 792 318
rect 838 272 870 318
rect 760 210 870 272
rect 930 318 1040 380
rect 930 272 962 318
rect 1008 272 1040 318
rect 930 210 1040 272
rect 1100 318 1210 380
rect 1100 272 1132 318
rect 1178 272 1210 318
rect 1100 210 1210 272
rect 1270 318 1380 380
rect 1270 272 1302 318
rect 1348 272 1380 318
rect 1270 210 1380 272
rect 1440 318 1550 380
rect 1440 272 1472 318
rect 1518 272 1550 318
rect 1440 210 1550 272
rect 1610 318 1720 380
rect 1610 272 1642 318
rect 1688 272 1720 318
rect 1610 210 1720 272
rect 1780 318 1890 380
rect 1780 272 1812 318
rect 1858 272 1890 318
rect 1780 210 1890 272
rect 1950 318 2060 380
rect 1950 272 1982 318
rect 2028 272 2060 318
rect 1950 210 2060 272
rect 2120 318 2230 380
rect 2120 272 2152 318
rect 2198 272 2230 318
rect 2120 210 2230 272
rect 2290 318 2400 380
rect 2290 272 2322 318
rect 2368 272 2400 318
rect 2290 210 2400 272
rect 2460 318 2570 380
rect 2460 272 2492 318
rect 2538 272 2570 318
rect 2460 210 2570 272
rect 2630 318 2740 380
rect 2630 272 2662 318
rect 2708 272 2740 318
rect 2630 210 2740 272
rect 2800 318 2910 380
rect 2800 272 2832 318
rect 2878 272 2910 318
rect 2800 210 2910 272
rect 2970 318 3070 380
rect 2970 272 3002 318
rect 3048 272 3070 318
rect 2970 210 3070 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1397 530 1450
rect 420 1163 452 1397
rect 498 1163 530 1397
rect 420 1110 530 1163
rect 590 1397 700 1450
rect 590 1163 622 1397
rect 668 1163 700 1397
rect 590 1110 700 1163
rect 760 1397 870 1450
rect 760 1163 792 1397
rect 838 1163 870 1397
rect 760 1110 870 1163
rect 930 1397 1040 1450
rect 930 1163 962 1397
rect 1008 1163 1040 1397
rect 930 1110 1040 1163
rect 1100 1397 1210 1450
rect 1100 1163 1132 1397
rect 1178 1163 1210 1397
rect 1100 1110 1210 1163
rect 1270 1397 1380 1450
rect 1270 1163 1302 1397
rect 1348 1163 1380 1397
rect 1270 1110 1380 1163
rect 1440 1397 1550 1450
rect 1440 1163 1472 1397
rect 1518 1163 1550 1397
rect 1440 1110 1550 1163
rect 1610 1397 1720 1450
rect 1610 1163 1642 1397
rect 1688 1163 1720 1397
rect 1610 1110 1720 1163
rect 1780 1397 1890 1450
rect 1780 1163 1812 1397
rect 1858 1163 1890 1397
rect 1780 1110 1890 1163
rect 1950 1397 2060 1450
rect 1950 1163 1982 1397
rect 2028 1163 2060 1397
rect 1950 1110 2060 1163
rect 2120 1397 2230 1450
rect 2120 1163 2152 1397
rect 2198 1163 2230 1397
rect 2120 1110 2230 1163
rect 2290 1397 2400 1450
rect 2290 1163 2322 1397
rect 2368 1163 2400 1397
rect 2290 1110 2400 1163
rect 2460 1397 2570 1450
rect 2460 1163 2492 1397
rect 2538 1163 2570 1397
rect 2460 1110 2570 1163
rect 2630 1397 2740 1450
rect 2630 1163 2662 1397
rect 2708 1163 2740 1397
rect 2630 1110 2740 1163
rect 2800 1397 2910 1450
rect 2800 1163 2832 1397
rect 2878 1163 2910 1397
rect 2800 1110 2910 1163
rect 2970 1397 3070 1450
rect 2970 1163 3002 1397
rect 3048 1163 3070 1397
rect 2970 1110 3070 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 792 272 838 318
rect 962 272 1008 318
rect 1132 272 1178 318
rect 1302 272 1348 318
rect 1472 272 1518 318
rect 1642 272 1688 318
rect 1812 272 1858 318
rect 1982 272 2028 318
rect 2152 272 2198 318
rect 2322 272 2368 318
rect 2492 272 2538 318
rect 2662 272 2708 318
rect 2832 272 2878 318
rect 3002 272 3048 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 452 1163 498 1397
rect 622 1163 668 1397
rect 792 1163 838 1397
rect 962 1163 1008 1397
rect 1132 1163 1178 1397
rect 1302 1163 1348 1397
rect 1472 1163 1518 1397
rect 1642 1163 1688 1397
rect 1812 1163 1858 1397
rect 1982 1163 2028 1397
rect 2152 1163 2198 1397
rect 2322 1163 2368 1397
rect 2492 1163 2538 1397
rect 2662 1163 2708 1397
rect 2832 1163 2878 1397
rect 3002 1163 3048 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
rect 2700 118 2850 140
rect 2700 72 2752 118
rect 2798 72 2850 118
rect 2700 50 2850 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1020 1588 1170 1610
rect 1020 1542 1072 1588
rect 1118 1542 1170 1588
rect 1020 1520 1170 1542
rect 1260 1588 1410 1610
rect 1260 1542 1312 1588
rect 1358 1542 1410 1588
rect 1260 1520 1410 1542
rect 1500 1588 1650 1610
rect 1500 1542 1552 1588
rect 1598 1542 1650 1588
rect 1500 1520 1650 1542
rect 1740 1588 1890 1610
rect 1740 1542 1792 1588
rect 1838 1542 1890 1588
rect 1740 1520 1890 1542
rect 1980 1588 2130 1610
rect 1980 1542 2032 1588
rect 2078 1542 2130 1588
rect 1980 1520 2130 1542
rect 2220 1588 2370 1610
rect 2220 1542 2272 1588
rect 2318 1542 2370 1588
rect 2220 1520 2370 1542
rect 2460 1588 2610 1610
rect 2460 1542 2512 1588
rect 2558 1542 2610 1588
rect 2460 1520 2610 1542
rect 2700 1588 2850 1610
rect 2700 1542 2752 1588
rect 2798 1542 2850 1588
rect 2700 1520 2850 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
rect 2752 72 2798 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1072 1542 1118 1588
rect 1312 1542 1358 1588
rect 1552 1542 1598 1588
rect 1792 1542 1838 1588
rect 2032 1542 2078 1588
rect 2272 1542 2318 1588
rect 2512 1542 2558 1588
rect 2752 1542 2798 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 530 1450 590 1500
rect 700 1450 760 1500
rect 870 1450 930 1500
rect 1040 1450 1100 1500
rect 1210 1450 1270 1500
rect 1380 1450 1440 1500
rect 1550 1450 1610 1500
rect 1720 1450 1780 1500
rect 1890 1450 1950 1500
rect 2060 1450 2120 1500
rect 2230 1450 2290 1500
rect 2400 1450 2460 1500
rect 2570 1450 2630 1500
rect 2740 1450 2800 1500
rect 2910 1450 2970 1500
rect 190 930 250 1110
rect 360 1090 420 1110
rect 530 1090 590 1110
rect 700 1090 760 1110
rect 870 1090 930 1110
rect 1040 1090 1100 1110
rect 1210 1090 1270 1110
rect 1380 1090 1440 1110
rect 1550 1090 1610 1110
rect 1720 1090 1780 1110
rect 1890 1090 1950 1110
rect 2060 1090 2120 1110
rect 2230 1090 2290 1110
rect 2400 1090 2460 1110
rect 2570 1090 2630 1110
rect 2740 1090 2800 1110
rect 2910 1090 2970 1110
rect 360 1030 2970 1090
rect 190 903 310 930
rect 190 857 237 903
rect 283 857 310 903
rect 190 830 310 857
rect 190 380 250 830
rect 360 690 420 1030
rect 300 653 420 690
rect 300 607 327 653
rect 373 607 420 653
rect 300 570 420 607
rect 360 460 420 570
rect 700 460 760 1030
rect 1040 460 1100 1030
rect 1380 460 1440 1030
rect 1720 460 1780 1030
rect 2060 460 2120 1030
rect 2400 460 2460 1030
rect 2740 460 2800 1030
rect 360 400 2970 460
rect 360 380 420 400
rect 530 380 590 400
rect 700 380 760 400
rect 870 380 930 400
rect 1040 380 1100 400
rect 1210 380 1270 400
rect 1380 380 1440 400
rect 1550 380 1610 400
rect 1720 380 1780 400
rect 1890 380 1950 400
rect 2060 380 2120 400
rect 2230 380 2290 400
rect 2400 380 2460 400
rect 2570 380 2630 400
rect 2740 380 2800 400
rect 2910 380 2970 400
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
rect 870 160 930 210
rect 1040 160 1100 210
rect 1210 160 1270 210
rect 1380 160 1440 210
rect 1550 160 1610 210
rect 1720 160 1780 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2400 160 2460 210
rect 2570 160 2630 210
rect 2740 160 2800 210
rect 2910 160 2970 210
<< polycontact >>
rect 237 857 283 903
rect 327 607 373 653
<< metal1 >>
rect 0 1588 3160 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1072 1588
rect 1118 1542 1312 1588
rect 1358 1542 1552 1588
rect 1598 1542 1792 1588
rect 1838 1542 2032 1588
rect 2078 1542 2272 1588
rect 2318 1542 2512 1588
rect 2558 1542 2752 1588
rect 2798 1542 3160 1588
rect 0 1520 3160 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 660 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 450 1397 500 1450
rect 450 1163 452 1397
rect 498 1163 500 1397
rect 450 1050 500 1163
rect 620 1397 670 1520
rect 620 1163 622 1397
rect 668 1163 670 1397
rect 620 1110 670 1163
rect 790 1397 840 1450
rect 790 1163 792 1397
rect 838 1163 840 1397
rect 790 1050 840 1163
rect 960 1397 1010 1520
rect 960 1163 962 1397
rect 1008 1163 1010 1397
rect 960 1110 1010 1163
rect 1130 1397 1180 1450
rect 1130 1163 1132 1397
rect 1178 1163 1180 1397
rect 1130 1050 1180 1163
rect 1300 1397 1350 1520
rect 1300 1163 1302 1397
rect 1348 1163 1350 1397
rect 1300 1110 1350 1163
rect 1470 1397 1520 1450
rect 1470 1163 1472 1397
rect 1518 1163 1520 1397
rect 1470 1050 1520 1163
rect 1640 1397 1690 1520
rect 1640 1163 1642 1397
rect 1688 1163 1690 1397
rect 1640 1110 1690 1163
rect 1810 1397 1860 1450
rect 1810 1163 1812 1397
rect 1858 1163 1860 1397
rect 1810 1050 1860 1163
rect 1980 1397 2030 1520
rect 1980 1163 1982 1397
rect 2028 1163 2030 1397
rect 1980 1110 2030 1163
rect 2150 1397 2200 1450
rect 2150 1163 2152 1397
rect 2198 1163 2200 1397
rect 2150 1050 2200 1163
rect 2320 1397 2370 1520
rect 2320 1163 2322 1397
rect 2368 1163 2370 1397
rect 2320 1110 2370 1163
rect 2490 1397 2540 1450
rect 2490 1163 2492 1397
rect 2538 1163 2540 1397
rect 2490 1050 2540 1163
rect 2660 1397 2710 1520
rect 2660 1163 2662 1397
rect 2708 1163 2710 1397
rect 2660 1110 2710 1163
rect 2830 1397 2880 1450
rect 2830 1163 2832 1397
rect 2878 1163 2880 1397
rect 2830 1050 2880 1163
rect 3000 1397 3050 1520
rect 3000 1163 3002 1397
rect 3048 1163 3050 1397
rect 3000 1110 3050 1163
rect 450 1046 2910 1050
rect 450 994 2834 1046
rect 2886 994 2910 1046
rect 450 990 2910 994
rect 210 906 310 910
rect 210 854 234 906
rect 286 854 310 906
rect 210 850 310 854
rect 110 653 400 660
rect 110 607 327 653
rect 373 607 400 653
rect 110 600 400 607
rect 110 318 160 600
rect 450 480 500 990
rect 790 480 840 990
rect 1130 480 1180 990
rect 1470 480 1520 990
rect 1810 480 1860 990
rect 2150 480 2200 990
rect 2490 480 2540 990
rect 2830 480 2880 990
rect 450 430 2880 480
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 450 318 500 430
rect 450 272 452 318
rect 498 272 500 318
rect 450 210 500 272
rect 620 318 670 380
rect 620 272 622 318
rect 668 272 670 318
rect 620 140 670 272
rect 790 318 840 430
rect 790 272 792 318
rect 838 272 840 318
rect 790 210 840 272
rect 960 318 1010 380
rect 960 272 962 318
rect 1008 272 1010 318
rect 960 140 1010 272
rect 1130 318 1180 430
rect 1130 272 1132 318
rect 1178 272 1180 318
rect 1130 210 1180 272
rect 1300 318 1350 380
rect 1300 272 1302 318
rect 1348 272 1350 318
rect 1300 140 1350 272
rect 1470 318 1520 430
rect 1470 272 1472 318
rect 1518 272 1520 318
rect 1470 210 1520 272
rect 1640 318 1690 380
rect 1640 272 1642 318
rect 1688 272 1690 318
rect 1640 140 1690 272
rect 1810 318 1860 430
rect 1810 272 1812 318
rect 1858 272 1860 318
rect 1810 210 1860 272
rect 1980 318 2030 380
rect 1980 272 1982 318
rect 2028 272 2030 318
rect 1980 140 2030 272
rect 2150 318 2200 430
rect 2150 272 2152 318
rect 2198 272 2200 318
rect 2150 210 2200 272
rect 2320 318 2370 380
rect 2320 272 2322 318
rect 2368 272 2370 318
rect 2320 140 2370 272
rect 2490 318 2540 430
rect 2490 272 2492 318
rect 2538 272 2540 318
rect 2490 210 2540 272
rect 2660 318 2710 380
rect 2660 272 2662 318
rect 2708 272 2710 318
rect 2660 140 2710 272
rect 2830 318 2880 430
rect 2830 272 2832 318
rect 2878 272 2880 318
rect 2830 210 2880 272
rect 3000 318 3050 380
rect 3000 272 3002 318
rect 3048 272 3050 318
rect 3000 140 3050 272
rect 0 118 3160 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2752 118
rect 2798 72 3160 118
rect 0 0 3160 72
<< via1 >>
rect 2834 994 2886 1046
rect 234 903 286 906
rect 234 857 237 903
rect 237 857 283 903
rect 283 857 286 903
rect 234 854 286 857
<< metal2 >>
rect 2810 1050 2910 1060
rect 2800 1046 2910 1050
rect 2800 994 2834 1046
rect 2886 994 2910 1046
rect 2800 990 2910 994
rect 2810 980 2910 990
rect 220 910 300 920
rect 210 906 310 910
rect 210 854 234 906
rect 286 854 310 906
rect 210 850 310 854
rect 220 840 300 850
<< labels >>
rlabel via1 s 234 854 286 906 4 A
port 1 nsew signal input
rlabel via1 s 2834 994 2886 1046 4 Y
port 2 nsew signal output
rlabel metal1 s 280 1110 330 1660 4 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 620 1110 670 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 960 1110 1010 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1300 1110 1350 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1640 1110 1690 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1980 1110 2030 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2320 1110 2370 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2660 1110 2710 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3000 1110 3050 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 1520 3160 1660 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 620 0 670 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 960 0 1010 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1300 0 1350 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1640 0 1690 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1980 0 2030 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2320 0 2370 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2660 0 2710 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3000 0 3050 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3160 140 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal2 s 220 840 300 920 1 A
port 1 nsew signal input
rlabel metal2 s 210 850 310 910 1 A
port 1 nsew signal input
rlabel metal1 s 210 850 310 910 1 A
port 1 nsew signal input
rlabel metal2 s 2800 990 2910 1050 1 Y
port 2 nsew signal output
rlabel metal2 s 2810 980 2910 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 450 210 500 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 790 210 840 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 1130 210 1180 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 1470 210 1520 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 1810 210 1860 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 2150 210 2200 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 2490 210 2540 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 450 430 2880 480 1 Y
port 2 nsew signal output
rlabel metal1 s 2830 210 2880 1450 1 Y
port 2 nsew signal output
rlabel metal1 s 450 990 2910 1050 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3160 1660
string GDS_END 133092
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 116292
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
