magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 758 1094
<< pwell >>
rect -86 -86 758 453
<< mvnmos >>
rect 124 187 244 333
rect 348 187 468 333
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
<< mvndiff >>
rect 36 246 124 333
rect 36 200 49 246
rect 95 200 124 246
rect 36 187 124 200
rect 244 246 348 333
rect 244 200 273 246
rect 319 200 348 246
rect 244 187 348 200
rect 468 246 556 333
rect 468 200 497 246
rect 543 200 556 246
rect 468 187 556 200
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 536 939
rect 448 721 477 861
rect 523 721 536 861
rect 448 573 536 721
<< mvndiffc >>
rect 49 200 95 246
rect 273 200 319 246
rect 497 200 543 246
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 124 513 224 573
rect 348 513 448 573
rect 70 500 448 513
rect 70 454 83 500
rect 317 454 448 500
rect 70 441 448 454
rect 124 333 244 441
rect 348 377 448 441
rect 348 333 468 377
rect 124 143 244 187
rect 348 143 468 187
<< polycontact >>
rect 83 454 317 500
<< metal1 >>
rect 0 918 672 1098
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 477 861 523 918
rect 319 721 420 766
rect 273 710 420 721
rect 477 710 523 721
rect 366 578 420 710
rect 72 500 328 542
rect 72 454 83 500
rect 317 454 328 500
rect 374 408 420 578
rect 273 362 420 408
rect 49 246 95 257
rect 49 90 95 200
rect 273 246 319 362
rect 273 189 319 200
rect 497 246 543 257
rect 497 90 543 200
rect 0 -90 672 90
<< labels >>
flabel metal1 s 72 454 328 542 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 672 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 497 90 543 257 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 273 766 319 872 0 FreeSans 200 0 0 0 ZN
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 273 710 420 766 1 ZN
port 2 nsew default output
rlabel metal1 s 366 578 420 710 1 ZN
port 2 nsew default output
rlabel metal1 s 374 408 420 578 1 ZN
port 2 nsew default output
rlabel metal1 s 273 362 420 408 1 ZN
port 2 nsew default output
rlabel metal1 s 273 189 319 362 1 ZN
port 2 nsew default output
rlabel metal1 s 477 710 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 90 95 257 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 672 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 1008
string GDS_END 1446214
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1443520
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
