magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1640 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
rect 870 210 930 380
rect 1040 210 1100 380
rect 1210 210 1270 380
rect 1380 210 1440 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
rect 700 720 760 1060
rect 870 720 930 1060
rect 1040 720 1100 1060
rect 1210 720 1270 1060
rect 1380 720 1440 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 318 530 380
rect 420 272 452 318
rect 498 272 530 318
rect 420 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 318 870 380
rect 760 272 792 318
rect 838 272 870 318
rect 760 210 870 272
rect 930 318 1040 380
rect 930 272 962 318
rect 1008 272 1040 318
rect 930 210 1040 272
rect 1100 318 1210 380
rect 1100 272 1132 318
rect 1178 272 1210 318
rect 1100 210 1210 272
rect 1270 318 1380 380
rect 1270 272 1302 318
rect 1348 272 1380 318
rect 1270 210 1380 272
rect 1440 318 1540 380
rect 1440 272 1472 318
rect 1518 272 1540 318
rect 1440 210 1540 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 360 1060
rect 250 773 282 1007
rect 328 773 360 1007
rect 250 720 360 773
rect 420 1007 530 1060
rect 420 773 452 1007
rect 498 773 530 1007
rect 420 720 530 773
rect 590 1007 700 1060
rect 590 773 622 1007
rect 668 773 700 1007
rect 590 720 700 773
rect 760 1007 870 1060
rect 760 773 792 1007
rect 838 773 870 1007
rect 760 720 870 773
rect 930 1007 1040 1060
rect 930 773 962 1007
rect 1008 773 1040 1007
rect 930 720 1040 773
rect 1100 1007 1210 1060
rect 1100 773 1132 1007
rect 1178 773 1210 1007
rect 1100 720 1210 773
rect 1270 1007 1380 1060
rect 1270 773 1302 1007
rect 1348 773 1380 1007
rect 1270 720 1380 773
rect 1440 1007 1550 1060
rect 1440 773 1482 1007
rect 1528 773 1550 1007
rect 1440 720 1550 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 792 272 838 318
rect 962 272 1008 318
rect 1132 272 1178 318
rect 1302 272 1348 318
rect 1472 272 1518 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 452 773 498 1007
rect 622 773 668 1007
rect 792 773 838 1007
rect 962 773 1008 1007
rect 1132 773 1178 1007
rect 1302 773 1348 1007
rect 1482 773 1528 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 700 1060 760 1110
rect 870 1060 930 1110
rect 1040 1060 1100 1110
rect 1210 1060 1270 1110
rect 1380 1060 1440 1110
rect 190 670 250 720
rect 360 670 420 720
rect 530 670 590 720
rect 700 670 760 720
rect 870 670 930 720
rect 1040 670 1100 720
rect 1210 670 1270 720
rect 1380 670 1440 720
rect 190 620 1440 670
rect 190 540 250 620
rect 90 518 250 540
rect 90 472 112 518
rect 158 480 250 518
rect 158 472 1440 480
rect 90 450 1440 472
rect 190 420 1440 450
rect 190 380 250 420
rect 360 380 420 420
rect 530 380 590 420
rect 700 380 760 420
rect 870 380 930 420
rect 1040 380 1100 420
rect 1210 380 1270 420
rect 1380 380 1440 420
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
rect 870 160 930 210
rect 1040 160 1100 210
rect 1210 160 1270 210
rect 1380 160 1440 210
<< polycontact >>
rect 112 472 158 518
<< metal1 >>
rect 0 1198 1640 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1640 1198
rect 0 1130 1640 1152
rect 110 1007 160 1130
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 720 160 773
rect 280 1007 330 1060
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 670 330 773
rect 450 1007 500 1130
rect 450 773 452 1007
rect 498 773 500 1007
rect 450 720 500 773
rect 620 1007 670 1060
rect 620 773 622 1007
rect 668 773 670 1007
rect 620 670 670 773
rect 790 1007 840 1130
rect 790 773 792 1007
rect 838 773 840 1007
rect 790 720 840 773
rect 960 1007 1010 1060
rect 960 773 962 1007
rect 1008 773 1010 1007
rect 960 670 1010 773
rect 1130 1007 1180 1130
rect 1130 773 1132 1007
rect 1178 773 1180 1007
rect 1130 720 1180 773
rect 1300 1007 1350 1060
rect 1300 773 1302 1007
rect 1348 780 1350 1007
rect 1480 1007 1530 1130
rect 1348 776 1430 780
rect 1348 773 1354 776
rect 1300 724 1354 773
rect 1406 724 1430 776
rect 1300 720 1430 724
rect 1480 773 1482 1007
rect 1528 773 1530 1007
rect 1480 720 1530 773
rect 1300 670 1350 720
rect 280 620 1350 670
rect 80 518 180 520
rect 80 516 112 518
rect 80 464 104 516
rect 158 472 180 518
rect 156 464 180 472
rect 80 460 180 464
rect 280 480 330 620
rect 620 480 670 620
rect 960 480 1010 620
rect 1300 480 1350 620
rect 280 430 1350 480
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 430
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 450 318 500 380
rect 450 272 452 318
rect 498 272 500 318
rect 450 140 500 272
rect 620 318 670 430
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 790 318 840 380
rect 790 272 792 318
rect 838 272 840 318
rect 790 140 840 272
rect 960 318 1010 430
rect 960 272 962 318
rect 1008 272 1010 318
rect 960 210 1010 272
rect 1130 318 1180 380
rect 1130 272 1132 318
rect 1178 272 1180 318
rect 1130 140 1180 272
rect 1300 318 1350 430
rect 1300 272 1302 318
rect 1348 272 1350 318
rect 1300 210 1350 272
rect 1470 318 1520 380
rect 1470 272 1472 318
rect 1518 272 1520 318
rect 1470 140 1520 272
rect 0 118 1640 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1640 118
rect 0 0 1640 72
<< via1 >>
rect 1354 724 1406 776
rect 104 472 112 516
rect 112 472 156 516
rect 104 464 156 472
<< metal2 >>
rect 1340 780 1420 790
rect 1330 776 1430 780
rect 1330 724 1354 776
rect 1406 724 1430 776
rect 1330 720 1430 724
rect 1340 710 1420 720
rect 80 516 180 530
rect 80 464 104 516
rect 156 464 180 516
rect 80 450 180 464
<< labels >>
rlabel via1 s 104 464 156 516 4 A
port 1 nsew signal input
rlabel via1 s 1354 724 1406 776 4 Y
port 2 nsew signal output
rlabel metal1 s 110 720 160 1270 4 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 110 0 160 380 4 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 450 720 500 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 790 720 840 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1130 720 1180 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1480 720 1530 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1640 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 450 0 500 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 790 0 840 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1130 0 1180 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1470 0 1520 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1640 140 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal2 s 80 450 180 530 1 A
port 1 nsew signal input
rlabel metal1 s 80 460 180 520 1 A
port 1 nsew signal input
rlabel metal2 s 1340 710 1420 790 1 Y
port 2 nsew signal output
rlabel metal2 s 1330 720 1430 780 1 Y
port 2 nsew signal output
rlabel metal1 s 280 210 330 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 620 210 670 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 960 210 1010 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 280 430 1350 480 1 Y
port 2 nsew signal output
rlabel metal1 s 280 620 1350 670 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 210 1350 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 720 1430 780 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1640 1270
string GDS_END 305540
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 296548
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
