magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 453 1990 1094
<< pwell >>
rect -86 -86 1990 453
<< mvnmos >>
rect 124 69 244 333
rect 396 201 516 333
rect 564 201 684 333
rect 932 201 1052 333
rect 1156 201 1276 333
rect 1380 201 1500 333
rect 1640 69 1760 333
<< mvpmos >>
rect 144 573 244 939
rect 396 691 496 874
rect 600 691 700 874
rect 952 691 1052 874
rect 1156 691 1256 874
rect 1400 691 1500 874
rect 1640 573 1740 939
<< mvndiff >>
rect 36 320 124 333
rect 36 180 49 320
rect 95 180 124 320
rect 36 69 124 180
rect 244 259 396 333
rect 244 213 273 259
rect 319 213 396 259
rect 244 201 396 213
rect 516 201 564 333
rect 684 260 772 333
rect 684 214 713 260
rect 759 214 772 260
rect 684 201 772 214
rect 844 260 932 333
rect 844 214 857 260
rect 903 214 932 260
rect 844 201 932 214
rect 1052 285 1156 333
rect 1052 239 1081 285
rect 1127 239 1156 285
rect 1052 201 1156 239
rect 1276 260 1380 333
rect 1276 214 1305 260
rect 1351 214 1380 260
rect 1276 201 1380 214
rect 1500 260 1640 333
rect 1500 214 1529 260
rect 1575 214 1640 260
rect 1500 201 1640 214
rect 244 69 324 201
rect 1560 69 1640 201
rect 1760 320 1848 333
rect 1760 180 1789 320
rect 1835 180 1848 320
rect 1760 69 1848 180
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 874 324 939
rect 1560 874 1640 939
rect 244 861 396 874
rect 244 721 273 861
rect 319 721 396 861
rect 244 691 396 721
rect 496 861 600 874
rect 496 721 525 861
rect 571 721 600 861
rect 496 691 600 721
rect 700 849 788 874
rect 700 803 729 849
rect 775 803 788 849
rect 700 691 788 803
rect 864 849 952 874
rect 864 803 877 849
rect 923 803 952 849
rect 864 691 952 803
rect 1052 691 1156 874
rect 1256 838 1400 874
rect 1256 792 1325 838
rect 1371 792 1400 838
rect 1256 691 1400 792
rect 1500 861 1640 874
rect 1500 721 1529 861
rect 1575 721 1640 861
rect 1500 691 1640 721
rect 244 573 324 691
rect 1560 573 1640 691
rect 1740 861 1828 939
rect 1740 721 1769 861
rect 1815 721 1828 861
rect 1740 573 1828 721
<< mvndiffc >>
rect 49 180 95 320
rect 273 213 319 259
rect 713 214 759 260
rect 857 214 903 260
rect 1081 239 1127 285
rect 1305 214 1351 260
rect 1529 214 1575 260
rect 1789 180 1835 320
<< mvpdiffc >>
rect 69 721 115 861
rect 273 721 319 861
rect 525 721 571 861
rect 729 803 775 849
rect 877 803 923 849
rect 1325 792 1371 838
rect 1529 721 1575 861
rect 1769 721 1815 861
<< polysilicon >>
rect 144 939 244 983
rect 1640 939 1740 983
rect 396 874 496 918
rect 600 874 700 918
rect 952 874 1052 918
rect 1156 874 1256 918
rect 1400 874 1500 918
rect 396 607 496 691
rect 396 594 516 607
rect 144 500 244 573
rect 144 454 185 500
rect 231 454 244 500
rect 144 377 244 454
rect 124 333 244 377
rect 396 454 457 594
rect 503 454 516 594
rect 600 513 700 691
rect 952 513 1052 691
rect 600 511 1052 513
rect 396 333 516 454
rect 564 500 1052 511
rect 564 454 607 500
rect 935 454 1052 500
rect 564 441 1052 454
rect 564 333 684 441
rect 932 333 1052 441
rect 1156 594 1256 691
rect 1156 454 1169 594
rect 1215 454 1256 594
rect 1156 377 1256 454
rect 1400 500 1500 691
rect 1400 454 1413 500
rect 1459 454 1500 500
rect 1400 377 1500 454
rect 1156 333 1276 377
rect 1380 333 1500 377
rect 1640 500 1740 573
rect 1640 454 1653 500
rect 1699 454 1740 500
rect 1640 377 1740 454
rect 1640 333 1760 377
rect 396 157 516 201
rect 564 157 684 201
rect 932 157 1052 201
rect 1156 157 1276 201
rect 1380 157 1500 201
rect 124 25 244 69
rect 1640 25 1760 69
<< polycontact >>
rect 185 454 231 500
rect 457 454 503 594
rect 607 454 935 500
rect 1169 454 1215 594
rect 1413 454 1459 500
rect 1653 454 1699 500
<< metal1 >>
rect 0 918 1904 1098
rect 30 861 115 872
rect 30 721 69 861
rect 30 320 115 721
rect 273 861 319 918
rect 525 861 571 872
rect 273 710 319 721
rect 365 721 525 746
rect 729 849 775 918
rect 729 792 775 803
rect 877 849 923 918
rect 1529 861 1575 918
rect 877 792 923 803
rect 1314 792 1325 838
rect 1371 792 1483 838
rect 571 721 1391 746
rect 365 700 1391 721
rect 365 511 411 700
rect 185 500 411 511
rect 231 454 411 500
rect 185 443 411 454
rect 457 594 1215 654
rect 503 590 1169 594
rect 590 500 1039 530
rect 590 454 607 500
rect 935 454 1039 500
rect 1345 500 1391 700
rect 1437 664 1483 792
rect 1529 710 1575 721
rect 1769 861 1835 872
rect 1815 721 1835 861
rect 1437 618 1562 664
rect 1516 511 1562 618
rect 1516 500 1699 511
rect 1345 454 1413 500
rect 1459 454 1470 500
rect 1516 454 1653 500
rect 457 443 503 454
rect 1169 443 1215 454
rect 1516 443 1699 454
rect 30 180 49 320
rect 95 180 115 320
rect 30 169 115 180
rect 273 259 319 270
rect 365 260 411 443
rect 1516 397 1562 443
rect 1081 351 1562 397
rect 1081 285 1127 351
rect 1769 320 1835 721
rect 1769 318 1789 320
rect 857 260 903 271
rect 365 214 713 260
rect 759 214 770 260
rect 1081 228 1127 239
rect 1305 260 1351 271
rect 273 90 319 213
rect 857 182 903 214
rect 1305 182 1351 214
rect 857 136 1351 182
rect 1529 260 1575 271
rect 1710 242 1789 318
rect 1529 90 1575 214
rect 1789 169 1835 180
rect 0 -90 1904 90
<< labels >>
flabel metal1 s 457 590 1215 654 0 FreeSans 200 0 0 0 A
port 1 nsew default input
flabel metal1 s 590 454 1039 530 0 FreeSans 200 0 0 0 B
port 2 nsew default input
flabel metal1 s 30 169 115 872 0 FreeSans 200 0 0 0 CO
port 3 nsew default output
flabel metal1 s 1769 318 1835 872 0 FreeSans 200 0 0 0 S
port 4 nsew default output
flabel metal1 s 0 918 1904 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1529 270 1575 271 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 1169 443 1215 590 1 A
port 1 nsew default input
rlabel metal1 s 457 443 503 590 1 A
port 1 nsew default input
rlabel metal1 s 1710 242 1835 318 1 S
port 4 nsew default output
rlabel metal1 s 1789 169 1835 242 1 S
port 4 nsew default output
rlabel metal1 s 1529 792 1575 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 877 792 923 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 729 792 775 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 792 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1529 710 1575 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 710 319 792 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1529 90 1575 270 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 270 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1904 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 1008
string GDS_END 1109168
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1103710
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
