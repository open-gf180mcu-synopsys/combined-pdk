magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 459 2326 1094
rect -86 453 86 459
rect 1871 453 2326 459
<< pwell >>
rect 86 453 1871 459
rect -86 -86 2326 453
<< mvnmos >>
rect 397 267 517 339
rect 124 123 244 195
rect 397 123 517 195
rect 829 212 949 284
rect 1197 212 1317 284
rect 829 68 949 140
rect 1197 68 1317 140
rect 1629 213 1749 285
rect 1629 69 1749 141
rect 1989 69 2109 333
<< mvpmos >>
rect 124 774 224 846
rect 397 774 497 846
rect 397 630 497 702
rect 829 774 929 846
rect 1197 774 1297 846
rect 829 630 929 702
rect 1197 630 1297 702
rect 1629 774 1729 846
rect 1629 630 1729 702
rect 1989 573 2089 939
<< mvndiff >>
rect 309 326 397 339
rect 309 280 322 326
rect 368 280 397 326
rect 309 267 397 280
rect 517 267 637 339
rect 577 195 637 267
rect 36 182 124 195
rect 36 136 49 182
rect 95 136 124 182
rect 36 123 124 136
rect 244 182 397 195
rect 244 136 273 182
rect 319 136 397 182
rect 244 123 397 136
rect 517 123 637 195
rect 709 212 829 284
rect 949 271 1037 284
rect 949 225 978 271
rect 1024 225 1037 271
rect 949 212 1037 225
rect 1109 271 1197 284
rect 1109 225 1122 271
rect 1168 225 1197 271
rect 1109 212 1197 225
rect 1317 212 1437 284
rect 709 140 769 212
rect 1377 140 1437 212
rect 709 68 829 140
rect 949 127 1197 140
rect 949 81 978 127
rect 1024 81 1197 127
rect 949 68 1197 81
rect 1317 68 1437 140
rect 1509 213 1629 285
rect 1749 272 1837 285
rect 1749 226 1778 272
rect 1824 226 1837 272
rect 1749 213 1837 226
rect 1509 141 1569 213
rect 1909 141 1989 333
rect 1509 69 1629 141
rect 1749 128 1989 141
rect 1749 82 1778 128
rect 1824 82 1989 128
rect 1749 69 1989 82
rect 2109 287 2197 333
rect 2109 147 2138 287
rect 2184 147 2197 287
rect 2109 69 2197 147
<< mvpdiff >>
rect 1909 846 1989 939
rect 36 833 124 846
rect 36 787 49 833
rect 95 787 124 833
rect 36 774 124 787
rect 224 833 397 846
rect 224 787 322 833
rect 368 787 397 833
rect 224 774 397 787
rect 497 774 617 846
rect 557 702 617 774
rect 309 689 397 702
rect 309 643 322 689
rect 368 643 397 689
rect 309 630 397 643
rect 497 630 617 702
rect 709 774 829 846
rect 929 833 1197 846
rect 929 787 958 833
rect 1004 787 1197 833
rect 929 774 1197 787
rect 1297 774 1417 846
rect 709 702 769 774
rect 1357 702 1417 774
rect 709 630 829 702
rect 929 689 1017 702
rect 929 643 958 689
rect 1004 643 1017 689
rect 929 630 1017 643
rect 1109 689 1197 702
rect 1109 643 1122 689
rect 1168 643 1197 689
rect 1109 630 1197 643
rect 1297 630 1417 702
rect 1509 774 1629 846
rect 1729 833 1989 846
rect 1729 787 1758 833
rect 1804 787 1989 833
rect 1729 774 1989 787
rect 1509 702 1569 774
rect 1509 630 1629 702
rect 1729 689 1817 702
rect 1729 643 1758 689
rect 1804 643 1817 689
rect 1729 630 1817 643
rect 1909 573 1989 774
rect 2089 861 2177 939
rect 2089 721 2118 861
rect 2164 721 2177 861
rect 2089 573 2177 721
<< mvndiffc >>
rect 322 280 368 326
rect 49 136 95 182
rect 273 136 319 182
rect 978 225 1024 271
rect 1122 225 1168 271
rect 978 81 1024 127
rect 1778 226 1824 272
rect 1778 82 1824 128
rect 2138 147 2184 287
<< mvpdiffc >>
rect 49 787 95 833
rect 322 787 368 833
rect 322 643 368 689
rect 958 787 1004 833
rect 958 643 1004 689
rect 1122 643 1168 689
rect 1758 787 1804 833
rect 1758 643 1804 689
rect 2118 721 2164 861
<< polysilicon >>
rect 1989 939 2089 983
rect 124 846 224 890
rect 397 846 497 890
rect 829 846 929 890
rect 1197 846 1297 890
rect 1629 846 1729 890
rect 124 512 224 774
rect 397 702 497 774
rect 829 702 929 774
rect 1197 702 1297 774
rect 1629 702 1729 774
rect 124 372 137 512
rect 183 372 224 512
rect 124 239 224 372
rect 397 512 497 630
rect 397 372 410 512
rect 456 383 497 512
rect 829 512 929 630
rect 456 372 517 383
rect 397 339 517 372
rect 829 372 842 512
rect 888 372 929 512
rect 829 328 929 372
rect 1197 512 1297 630
rect 1197 372 1210 512
rect 1256 372 1297 512
rect 1197 328 1297 372
rect 1629 512 1729 630
rect 1629 372 1642 512
rect 1688 372 1729 512
rect 1629 329 1729 372
rect 1989 512 2089 573
rect 1989 372 2002 512
rect 2048 377 2089 512
rect 2048 372 2109 377
rect 1989 333 2109 372
rect 829 284 949 328
rect 1197 284 1317 328
rect 1629 285 1749 329
rect 124 195 244 239
rect 397 195 517 267
rect 829 140 949 212
rect 1197 140 1317 212
rect 124 79 244 123
rect 397 79 517 123
rect 1629 141 1749 213
rect 829 24 949 68
rect 1197 24 1317 68
rect 1629 25 1749 69
rect 1989 25 2109 69
<< polycontact >>
rect 137 372 183 512
rect 410 372 456 512
rect 842 372 888 512
rect 1210 372 1256 512
rect 1642 372 1688 512
rect 2002 372 2048 512
<< metal1 >>
rect 0 918 2240 1098
rect 322 844 368 918
rect 2118 861 2184 872
rect 34 833 95 844
rect 34 787 49 833
rect 34 604 95 787
rect 322 833 1804 844
rect 368 787 958 833
rect 1004 787 1758 833
rect 322 776 1804 787
rect 2164 721 2184 861
rect 958 689 1004 700
rect 311 643 322 689
rect 368 643 888 689
rect 34 558 286 604
rect 34 182 80 558
rect 240 512 286 558
rect 842 512 888 643
rect 126 372 137 512
rect 183 372 194 512
rect 240 466 410 512
rect 399 372 410 466
rect 456 372 467 512
rect 126 354 194 372
rect 842 326 888 372
rect 311 280 322 326
rect 368 280 888 326
rect 958 418 1004 643
rect 1122 689 1168 700
rect 1122 604 1168 643
rect 1758 689 1804 700
rect 2118 654 2184 721
rect 1122 558 1359 604
rect 1199 418 1210 512
rect 958 372 1210 418
rect 1256 372 1267 512
rect 958 271 1024 372
rect 1313 326 1359 558
rect 1642 512 1688 523
rect 1642 326 1688 372
rect 958 225 978 271
rect 958 214 1024 225
rect 1122 280 1688 326
rect 1758 418 1804 643
rect 2046 578 2184 654
rect 1991 418 2002 512
rect 1758 372 2002 418
rect 2048 372 2059 512
rect 1122 271 1168 280
rect 1122 214 1168 225
rect 1758 272 1824 372
rect 1758 226 1778 272
rect 1758 215 1824 226
rect 2138 287 2184 578
rect 273 182 319 193
rect 34 136 49 182
rect 95 136 106 182
rect 273 90 319 136
rect 978 127 1024 138
rect 0 81 978 90
rect 1778 128 1824 139
rect 2138 136 2184 147
rect 1024 82 1778 90
rect 1824 82 2240 90
rect 1024 81 2240 82
rect 0 -90 2240 81
<< labels >>
flabel metal1 s 126 354 194 512 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 2240 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 273 139 319 193 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2118 654 2184 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2046 578 2184 654 1 Z
port 2 nsew default output
rlabel metal1 s 2138 136 2184 578 1 Z
port 2 nsew default output
rlabel metal1 s 322 844 368 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 322 776 1804 844 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1778 138 1824 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 138 319 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1778 90 1824 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 978 90 1024 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2240 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2240 1008
string GDS_END 727580
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 722070
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
