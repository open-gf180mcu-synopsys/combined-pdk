magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 2800 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
rect 870 210 930 380
rect 1040 210 1100 380
rect 1210 210 1270 380
rect 1380 210 1440 380
rect 1550 210 1610 380
rect 1720 210 1780 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2550 210 2610 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
rect 700 720 760 1060
rect 870 720 930 1060
rect 1040 720 1100 1060
rect 1210 720 1270 1060
rect 1380 720 1440 1060
rect 1550 720 1610 1060
rect 1720 720 1780 1060
rect 1890 720 1950 1060
rect 2060 720 2120 1060
rect 2230 720 2290 1060
rect 2550 720 2610 1060
<< ndiff >>
rect 90 278 190 380
rect 90 232 112 278
rect 158 232 190 278
rect 90 210 190 232
rect 250 278 360 380
rect 250 232 282 278
rect 328 232 360 278
rect 250 210 360 232
rect 420 278 530 380
rect 420 232 452 278
rect 498 232 530 278
rect 420 210 530 232
rect 590 278 700 380
rect 590 232 622 278
rect 668 232 700 278
rect 590 210 700 232
rect 760 210 870 380
rect 930 278 1040 380
rect 930 232 962 278
rect 1008 232 1040 278
rect 930 210 1040 232
rect 1100 278 1210 380
rect 1100 232 1132 278
rect 1178 232 1210 278
rect 1100 210 1210 232
rect 1270 278 1380 380
rect 1270 232 1302 278
rect 1348 232 1380 278
rect 1270 210 1380 232
rect 1440 278 1550 380
rect 1440 232 1472 278
rect 1518 232 1550 278
rect 1440 210 1550 232
rect 1610 278 1720 380
rect 1610 232 1642 278
rect 1688 232 1720 278
rect 1610 210 1720 232
rect 1780 210 1890 380
rect 1950 210 2060 380
rect 2120 278 2230 380
rect 2120 232 2152 278
rect 2198 232 2230 278
rect 2120 210 2230 232
rect 2290 278 2390 380
rect 2290 232 2322 278
rect 2368 232 2390 278
rect 2290 210 2390 232
rect 2450 278 2550 380
rect 2450 232 2472 278
rect 2518 232 2550 278
rect 2450 210 2550 232
rect 2610 278 2710 380
rect 2610 232 2642 278
rect 2688 232 2710 278
rect 2610 210 2710 232
<< pdiff >>
rect 90 1033 190 1060
rect 90 987 112 1033
rect 158 987 190 1033
rect 90 720 190 987
rect 250 1033 360 1060
rect 250 987 282 1033
rect 328 987 360 1033
rect 250 720 360 987
rect 420 1033 530 1060
rect 420 987 452 1033
rect 498 987 530 1033
rect 420 720 530 987
rect 590 1038 700 1060
rect 590 992 622 1038
rect 668 992 700 1038
rect 590 720 700 992
rect 760 720 870 1060
rect 930 1033 1040 1060
rect 930 987 962 1033
rect 1008 987 1040 1033
rect 930 720 1040 987
rect 1100 1033 1210 1060
rect 1100 987 1132 1033
rect 1178 987 1210 1033
rect 1100 720 1210 987
rect 1270 1033 1380 1060
rect 1270 987 1302 1033
rect 1348 987 1380 1033
rect 1270 720 1380 987
rect 1440 1033 1550 1060
rect 1440 987 1472 1033
rect 1518 987 1550 1033
rect 1440 720 1550 987
rect 1610 903 1720 1060
rect 1610 857 1642 903
rect 1688 857 1720 903
rect 1610 720 1720 857
rect 1780 720 1890 1060
rect 1950 720 2060 1060
rect 2120 1033 2230 1060
rect 2120 987 2152 1033
rect 2198 987 2230 1033
rect 2120 720 2230 987
rect 2290 1033 2390 1060
rect 2290 987 2322 1033
rect 2368 987 2390 1033
rect 2290 720 2390 987
rect 2450 1033 2550 1060
rect 2450 987 2472 1033
rect 2518 987 2550 1033
rect 2450 720 2550 987
rect 2610 1033 2710 1060
rect 2610 987 2642 1033
rect 2688 987 2710 1033
rect 2610 720 2710 987
<< ndiffc >>
rect 112 232 158 278
rect 282 232 328 278
rect 452 232 498 278
rect 622 232 668 278
rect 962 232 1008 278
rect 1132 232 1178 278
rect 1302 232 1348 278
rect 1472 232 1518 278
rect 1642 232 1688 278
rect 2152 232 2198 278
rect 2322 232 2368 278
rect 2472 232 2518 278
rect 2642 232 2688 278
<< pdiffc >>
rect 112 987 158 1033
rect 282 987 328 1033
rect 452 987 498 1033
rect 622 992 668 1038
rect 962 987 1008 1033
rect 1132 987 1178 1033
rect 1302 987 1348 1033
rect 1472 987 1518 1033
rect 1642 857 1688 903
rect 2152 987 2198 1033
rect 2322 987 2368 1033
rect 2472 987 2518 1033
rect 2642 987 2688 1033
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
rect 1500 1198 1650 1220
rect 1500 1152 1552 1198
rect 1598 1152 1650 1198
rect 1500 1130 1650 1152
rect 1740 1198 1890 1220
rect 1740 1152 1792 1198
rect 1838 1152 1890 1198
rect 1740 1130 1890 1152
rect 1980 1198 2130 1220
rect 1980 1152 2032 1198
rect 2078 1152 2130 1198
rect 1980 1130 2130 1152
rect 2220 1198 2370 1220
rect 2220 1152 2272 1198
rect 2318 1152 2370 1198
rect 2220 1130 2370 1152
rect 2460 1198 2610 1220
rect 2460 1152 2512 1198
rect 2558 1152 2610 1198
rect 2460 1130 2610 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
rect 1552 1152 1598 1198
rect 1792 1152 1838 1198
rect 2032 1152 2078 1198
rect 2272 1152 2318 1198
rect 2512 1152 2558 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 700 1060 760 1110
rect 870 1060 930 1110
rect 1040 1060 1100 1110
rect 1210 1060 1270 1110
rect 1380 1060 1440 1110
rect 1550 1060 1610 1110
rect 1720 1060 1780 1110
rect 1890 1060 1950 1110
rect 2060 1060 2120 1110
rect 2230 1060 2290 1110
rect 2550 1060 2610 1110
rect 190 540 250 720
rect 360 670 420 720
rect 300 643 420 670
rect 300 597 327 643
rect 373 597 420 643
rect 300 570 420 597
rect 120 513 250 540
rect 120 467 147 513
rect 193 467 250 513
rect 120 440 250 467
rect 190 380 250 440
rect 360 380 420 570
rect 530 540 590 720
rect 700 700 760 720
rect 870 700 930 720
rect 1040 700 1100 720
rect 1210 700 1270 720
rect 700 673 820 700
rect 700 627 747 673
rect 793 627 820 673
rect 700 600 820 627
rect 870 650 1100 700
rect 1150 673 1270 700
rect 510 513 610 540
rect 510 467 537 513
rect 583 467 610 513
rect 510 440 610 467
rect 530 380 590 440
rect 700 380 760 600
rect 870 570 930 650
rect 1150 627 1177 673
rect 1223 627 1270 673
rect 1150 600 1270 627
rect 870 543 1020 570
rect 870 497 947 543
rect 993 497 1020 543
rect 870 470 1020 497
rect 870 420 1100 470
rect 870 380 930 420
rect 1040 380 1100 420
rect 1210 380 1270 600
rect 1380 570 1440 720
rect 1550 570 1610 720
rect 1720 570 1780 720
rect 1890 700 1950 720
rect 1890 673 2010 700
rect 1890 627 1937 673
rect 1983 627 2010 673
rect 1890 600 2010 627
rect 1380 543 1490 570
rect 1380 497 1417 543
rect 1463 497 1490 543
rect 1380 470 1490 497
rect 1550 543 1660 570
rect 1550 497 1587 543
rect 1633 497 1660 543
rect 1550 470 1660 497
rect 1720 543 1840 570
rect 1720 497 1767 543
rect 1813 497 1840 543
rect 1720 470 1840 497
rect 1380 380 1440 470
rect 1550 380 1610 470
rect 1720 380 1780 470
rect 1890 380 1950 600
rect 2060 550 2120 720
rect 2230 570 2290 720
rect 2550 570 2610 720
rect 2020 523 2120 550
rect 2020 477 2047 523
rect 2093 477 2120 523
rect 2020 450 2120 477
rect 2170 543 2290 570
rect 2170 497 2197 543
rect 2243 497 2290 543
rect 2170 470 2290 497
rect 2490 543 2610 570
rect 2490 497 2517 543
rect 2563 497 2610 543
rect 2490 470 2610 497
rect 2060 380 2120 450
rect 2230 380 2290 470
rect 2550 380 2610 470
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
rect 870 160 930 210
rect 1040 160 1100 210
rect 1210 160 1270 210
rect 1380 160 1440 210
rect 1550 160 1610 210
rect 1720 160 1780 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2550 160 2610 210
<< polycontact >>
rect 327 597 373 643
rect 147 467 193 513
rect 747 627 793 673
rect 537 467 583 513
rect 1177 627 1223 673
rect 947 497 993 543
rect 1937 627 1983 673
rect 1417 497 1463 543
rect 1587 497 1633 543
rect 1767 497 1813 543
rect 2047 477 2093 523
rect 2197 497 2243 543
rect 2517 497 2563 543
<< metal1 >>
rect 0 1198 2800 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1552 1198
rect 1598 1152 1792 1198
rect 1838 1152 2032 1198
rect 2078 1152 2272 1198
rect 2318 1152 2512 1198
rect 2558 1152 2800 1198
rect 0 1130 2800 1152
rect 110 1033 160 1060
rect 110 987 112 1033
rect 158 987 160 1033
rect 110 910 160 987
rect 280 1033 330 1130
rect 280 987 282 1033
rect 328 987 330 1033
rect 280 960 330 987
rect 450 1033 500 1060
rect 450 987 452 1033
rect 498 987 500 1033
rect 450 910 500 987
rect 620 1038 680 1060
rect 620 992 622 1038
rect 668 1036 680 1038
rect 620 984 624 992
rect 676 984 680 1036
rect 620 960 680 984
rect 960 1033 1010 1130
rect 960 987 962 1033
rect 1008 987 1010 1033
rect 960 960 1010 987
rect 1130 1033 1180 1060
rect 1130 987 1132 1033
rect 1178 987 1180 1033
rect 110 860 500 910
rect 1130 910 1180 987
rect 1300 1033 1350 1130
rect 1300 987 1302 1033
rect 1348 987 1350 1033
rect 1300 960 1350 987
rect 1470 1033 1520 1060
rect 1470 987 1472 1033
rect 1518 987 1520 1033
rect 1470 910 1520 987
rect 2150 1033 2200 1130
rect 2150 987 2152 1033
rect 2198 987 2200 1033
rect 2150 960 2200 987
rect 2320 1033 2370 1060
rect 2320 987 2322 1033
rect 2368 987 2370 1033
rect 1130 860 1520 910
rect 1620 906 1720 910
rect 1620 903 1644 906
rect 1620 857 1642 903
rect 1620 854 1644 857
rect 1696 854 1720 906
rect 1620 850 1720 854
rect 320 750 800 810
rect 320 646 380 750
rect 320 594 324 646
rect 376 594 380 646
rect 320 570 380 594
rect 430 640 690 700
rect 430 520 480 640
rect 640 550 690 640
rect 740 680 800 750
rect 1170 740 1990 800
rect 1170 680 1230 740
rect 740 673 1230 680
rect 740 627 747 673
rect 793 627 1177 673
rect 1223 627 1230 673
rect 740 620 1230 627
rect 740 600 800 620
rect 1170 600 1230 620
rect 1280 630 1820 690
rect 1280 550 1340 630
rect 640 543 1340 550
rect 120 516 480 520
rect 120 464 144 516
rect 196 464 480 516
rect 120 460 480 464
rect 530 516 590 540
rect 530 464 534 516
rect 586 464 590 516
rect 640 497 947 543
rect 993 497 1340 543
rect 640 490 1340 497
rect 1410 543 1470 570
rect 1760 550 1820 630
rect 1930 673 1990 740
rect 1930 627 1937 673
rect 1983 627 1990 673
rect 1930 600 1990 627
rect 2320 690 2370 987
rect 2470 1033 2520 1130
rect 2470 987 2472 1033
rect 2518 987 2520 1033
rect 2470 960 2520 987
rect 2640 1033 2690 1060
rect 2640 987 2642 1033
rect 2688 987 2690 1033
rect 2640 690 2690 987
rect 2320 680 2380 690
rect 2640 680 2730 690
rect 2320 676 2410 680
rect 2320 624 2334 676
rect 2386 624 2410 676
rect 2320 620 2410 624
rect 2640 676 2750 680
rect 2640 624 2674 676
rect 2726 624 2750 676
rect 2640 620 2750 624
rect 2320 610 2380 620
rect 2640 610 2730 620
rect 1410 497 1417 543
rect 1463 497 1470 543
rect 530 440 590 464
rect 1410 440 1470 497
rect 1560 546 1660 550
rect 1560 494 1584 546
rect 1636 494 1660 546
rect 1560 490 1660 494
rect 1740 543 1840 550
rect 1740 497 1767 543
rect 1813 497 1840 543
rect 2170 546 2270 550
rect 1740 490 1840 497
rect 1950 523 2120 530
rect 1950 477 2047 523
rect 2093 477 2120 523
rect 2170 494 2194 546
rect 2246 494 2270 546
rect 2170 490 2270 494
rect 1950 470 2120 477
rect 1950 440 2010 470
rect 530 380 2010 440
rect 100 286 160 310
rect 100 234 104 286
rect 156 278 160 286
rect 100 232 112 234
rect 158 232 160 278
rect 100 210 160 232
rect 280 278 330 300
rect 280 232 282 278
rect 328 232 330 278
rect 280 140 330 232
rect 440 286 500 310
rect 440 234 444 286
rect 496 278 500 286
rect 440 232 452 234
rect 498 232 500 278
rect 440 210 500 232
rect 620 286 680 310
rect 620 278 624 286
rect 620 232 622 278
rect 676 234 680 286
rect 668 232 680 234
rect 620 210 680 232
rect 960 278 1010 300
rect 960 232 962 278
rect 1008 232 1010 278
rect 960 140 1010 232
rect 1130 286 1190 310
rect 1130 278 1134 286
rect 1130 232 1132 278
rect 1186 234 1190 286
rect 1178 232 1190 234
rect 1130 210 1190 232
rect 1300 278 1350 300
rect 1300 232 1302 278
rect 1348 232 1350 278
rect 1300 140 1350 232
rect 1460 286 1520 310
rect 1460 234 1464 286
rect 1516 278 1520 286
rect 1460 232 1472 234
rect 1518 232 1520 278
rect 1460 210 1520 232
rect 1640 286 1700 310
rect 1640 278 1644 286
rect 1640 232 1642 278
rect 1696 234 1700 286
rect 1688 232 1700 234
rect 1640 210 1700 232
rect 2150 278 2200 300
rect 2150 232 2152 278
rect 2198 232 2200 278
rect 2150 140 2200 232
rect 2320 278 2370 610
rect 2490 546 2590 550
rect 2490 494 2514 546
rect 2566 494 2590 546
rect 2490 490 2590 494
rect 2320 232 2322 278
rect 2368 232 2370 278
rect 2320 210 2370 232
rect 2470 278 2520 300
rect 2470 232 2472 278
rect 2518 232 2520 278
rect 2470 140 2520 232
rect 2640 278 2690 610
rect 2640 232 2642 278
rect 2688 232 2690 278
rect 2640 210 2690 232
rect 0 118 2800 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2800 118
rect 0 0 2800 72
<< via1 >>
rect 624 992 668 1036
rect 668 992 676 1036
rect 624 984 676 992
rect 1644 903 1696 906
rect 1644 857 1688 903
rect 1688 857 1696 903
rect 1644 854 1696 857
rect 324 643 376 646
rect 324 597 327 643
rect 327 597 373 643
rect 373 597 376 643
rect 324 594 376 597
rect 144 513 196 516
rect 144 467 147 513
rect 147 467 193 513
rect 193 467 196 513
rect 144 464 196 467
rect 534 513 586 516
rect 534 467 537 513
rect 537 467 583 513
rect 583 467 586 513
rect 534 464 586 467
rect 2334 624 2386 676
rect 2674 624 2726 676
rect 1584 543 1636 546
rect 1584 497 1587 543
rect 1587 497 1633 543
rect 1633 497 1636 543
rect 1584 494 1636 497
rect 2194 543 2246 546
rect 2194 497 2197 543
rect 2197 497 2243 543
rect 2243 497 2246 543
rect 2194 494 2246 497
rect 104 278 156 286
rect 104 234 112 278
rect 112 234 156 278
rect 444 278 496 286
rect 444 234 452 278
rect 452 234 496 278
rect 624 278 676 286
rect 624 234 668 278
rect 668 234 676 278
rect 1134 278 1186 286
rect 1134 234 1178 278
rect 1178 234 1186 278
rect 1464 278 1516 286
rect 1464 234 1472 278
rect 1472 234 1516 278
rect 1644 278 1696 286
rect 1644 234 1688 278
rect 1688 234 1696 278
rect 2514 543 2566 546
rect 2514 497 2517 543
rect 2517 497 2563 543
rect 2563 497 2566 543
rect 2514 494 2566 497
<< metal2 >>
rect 620 1050 680 1060
rect 610 1040 690 1050
rect 600 1036 2570 1040
rect 600 984 624 1036
rect 676 984 2570 1036
rect 600 980 2570 984
rect 610 970 690 980
rect 310 650 390 660
rect 300 646 400 650
rect 300 594 324 646
rect 376 594 400 646
rect 300 590 400 594
rect 310 580 390 590
rect 750 550 810 980
rect 1630 910 1710 920
rect 1620 906 2250 910
rect 1620 854 1644 906
rect 1696 854 2250 906
rect 1620 850 2250 854
rect 1630 840 1710 850
rect 1570 550 1650 560
rect 750 546 1660 550
rect 120 516 220 530
rect 520 520 600 530
rect 120 464 144 516
rect 196 464 220 516
rect 120 450 220 464
rect 510 516 610 520
rect 510 464 534 516
rect 586 464 610 516
rect 510 460 610 464
rect 750 494 1584 546
rect 1636 494 1660 546
rect 750 490 1660 494
rect 520 450 600 460
rect 100 300 160 310
rect 440 300 500 310
rect 620 300 680 310
rect 90 290 170 300
rect 430 290 510 300
rect 90 286 510 290
rect 90 234 104 286
rect 156 234 444 286
rect 496 234 510 286
rect 90 230 510 234
rect 90 220 170 230
rect 430 220 510 230
rect 610 290 690 300
rect 750 290 810 490
rect 1570 480 1650 490
rect 1130 300 1190 310
rect 1460 300 1520 310
rect 610 286 810 290
rect 610 234 624 286
rect 676 234 810 286
rect 610 230 810 234
rect 1120 290 1200 300
rect 1450 290 1530 300
rect 1630 290 1710 300
rect 1770 290 1830 850
rect 2190 560 2250 850
rect 2320 680 2400 690
rect 2310 676 2410 680
rect 2310 624 2334 676
rect 2386 624 2410 676
rect 2310 620 2410 624
rect 2320 610 2400 620
rect 2510 560 2570 980
rect 2660 680 2740 690
rect 2650 676 2750 680
rect 2650 624 2674 676
rect 2726 624 2750 676
rect 2650 620 2750 624
rect 2660 610 2740 620
rect 2180 546 2260 560
rect 2500 550 2580 560
rect 2180 494 2194 546
rect 2246 494 2260 546
rect 2180 480 2260 494
rect 2490 546 2590 550
rect 2490 494 2514 546
rect 2566 494 2590 546
rect 2490 490 2590 494
rect 2500 480 2580 490
rect 2190 470 2250 480
rect 2510 470 2570 480
rect 1120 286 1530 290
rect 1120 234 1134 286
rect 1186 234 1464 286
rect 1516 234 1530 286
rect 1120 230 1530 234
rect 1620 286 1830 290
rect 1620 234 1644 286
rect 1696 234 1830 286
rect 1620 230 1830 234
rect 610 220 690 230
rect 1120 220 1200 230
rect 1450 220 1530 230
rect 1630 220 1710 230
rect 100 210 160 220
rect 440 210 500 220
rect 620 210 680 220
rect 1130 210 1190 220
rect 1460 210 1520 220
<< labels >>
rlabel via1 s 144 464 196 516 4 A
port 1 nsew signal input
rlabel via1 s 324 594 376 646 4 B
port 2 nsew signal input
rlabel via1 s 534 464 586 516 4 CI
port 3 nsew signal input
rlabel via1 s 2334 624 2386 676 4 S
port 4 nsew signal output
rlabel via1 s 2674 624 2726 676 4 CO
port 5 nsew signal output
rlabel metal1 s 280 960 330 1270 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 300 4 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 960 960 1010 1270 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1300 960 1350 1270 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 960 2200 1270 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2470 960 2520 1270 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1130 2800 1270 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 960 0 1010 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1300 0 1350 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2150 0 2200 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2470 0 2520 300 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 0 2800 140 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal2 s 120 450 220 530 1 A
port 1 nsew signal input
rlabel metal1 s 120 460 480 520 1 A
port 1 nsew signal input
rlabel metal1 s 430 460 480 700 1 A
port 1 nsew signal input
rlabel metal1 s 640 490 690 700 1 A
port 1 nsew signal input
rlabel metal1 s 430 640 690 700 1 A
port 1 nsew signal input
rlabel metal1 s 640 490 1340 550 1 A
port 1 nsew signal input
rlabel metal1 s 1280 490 1340 690 1 A
port 1 nsew signal input
rlabel metal1 s 1760 490 1820 690 1 A
port 1 nsew signal input
rlabel metal1 s 1280 630 1820 690 1 A
port 1 nsew signal input
rlabel metal1 s 1740 490 1840 550 1 A
port 1 nsew signal input
rlabel metal2 s 310 580 390 660 1 B
port 2 nsew signal input
rlabel metal2 s 300 590 400 650 1 B
port 2 nsew signal input
rlabel metal1 s 320 570 380 810 1 B
port 2 nsew signal input
rlabel metal1 s 740 600 800 810 1 B
port 2 nsew signal input
rlabel metal1 s 320 750 800 810 1 B
port 2 nsew signal input
rlabel metal1 s 740 620 1230 680 1 B
port 2 nsew signal input
rlabel metal1 s 1170 600 1230 800 1 B
port 2 nsew signal input
rlabel metal1 s 1930 600 1990 800 1 B
port 2 nsew signal input
rlabel metal1 s 1170 740 1990 800 1 B
port 2 nsew signal input
rlabel metal2 s 520 450 600 530 1 CI
port 3 nsew signal input
rlabel metal2 s 510 460 610 520 1 CI
port 3 nsew signal input
rlabel metal1 s 530 380 590 540 1 CI
port 3 nsew signal input
rlabel metal1 s 1410 380 1470 570 1 CI
port 3 nsew signal input
rlabel metal1 s 530 380 2010 440 1 CI
port 3 nsew signal input
rlabel metal1 s 1950 380 2010 530 1 CI
port 3 nsew signal input
rlabel metal1 s 1950 470 2120 530 1 CI
port 3 nsew signal input
rlabel metal2 s 2660 610 2740 690 1 CO
port 5 nsew signal output
rlabel metal2 s 2650 620 2750 680 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 210 2690 1060 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 610 2730 690 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 620 2750 680 1 CO
port 5 nsew signal output
rlabel metal2 s 2320 610 2400 690 1 S
port 4 nsew signal output
rlabel metal2 s 2310 620 2410 680 1 S
port 4 nsew signal output
rlabel metal1 s 2320 210 2370 1060 1 S
port 4 nsew signal output
rlabel metal1 s 2320 610 2380 690 1 S
port 4 nsew signal output
rlabel metal1 s 2320 620 2410 680 1 S
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2800 1270
string GDS_END 19748
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 146
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
