VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__bi_24t
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_fd_io__bi_24t ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 264.310 69.780 350.000 ;
    END
  END A
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 328.395 3.740 350.000 ;
    END
  END CS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 72.435 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 55.175 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 23.680 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 17.930 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 9.070 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 17.930 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 17.930 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 9.815 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 2.320 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 9.040 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 9.040 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 9.040 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 9.040 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 2.310 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 60.835 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 60.835 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 60.835 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 71.955 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 66.365 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 59.650 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 52.120 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 54.080 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 63.560 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 68.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 9.320 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 9.320 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 19.780 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 19.735 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 2.985 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
  END DVSS
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.385 334.770 11.765 350.000 ;
    END
  END IE
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 7.776000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 266.190 70.510 350.000 ;
    END
  END OE
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 335.279999 ;
    PORT
      LAYER Metal3 ;
        RECT 25.000 20.000 50.000 45.000 ;
    END
  END PAD
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.330 329.950 10.710 350.000 ;
    END
  END PD
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.350000 ;
    ANTENNADIFFAREA 2.980000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.965 330.270 6.345 350.000 ;
    END
  END PU
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.670 264.990 69.050 350.000 ;
    END
  END SL
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 56.170 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 71.290 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.800000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.860 319.750 71.240 350.000 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 328.095 3.060 348.225 ;
        RECT 4.040 329.970 5.665 348.225 ;
        RECT 6.645 329.970 10.030 348.225 ;
        RECT 4.040 329.650 10.030 329.970 ;
        RECT 11.010 334.470 11.085 348.225 ;
        RECT 12.065 334.470 68.370 348.225 ;
        RECT 11.010 329.650 68.370 334.470 ;
        RECT 4.040 328.095 68.370 329.650 ;
        RECT 0.000 264.690 68.370 328.095 ;
        RECT 71.540 319.450 75.000 348.225 ;
        RECT 70.810 265.890 75.000 319.450 ;
        RECT 0.000 264.010 69.100 264.690 ;
        RECT 70.080 264.010 75.000 265.890 ;
        RECT 0.000 0.000 75.000 264.010 ;
      LAYER Metal3 ;
        RECT 11.120 342.800 66.200 348.390 ;
        RECT 25.480 340.200 66.200 342.800 ;
        RECT 25.480 334.800 71.790 340.200 ;
        RECT 25.480 332.200 61.760 334.800 ;
        RECT 11.120 324.200 61.760 332.200 ;
        RECT 2.800 318.800 72.200 324.200 ;
        RECT 2.800 310.800 69.490 318.800 ;
        RECT 21.580 300.200 52.280 310.800 ;
        RECT 19.730 294.800 53.375 300.200 ;
        RECT 21.535 284.200 50.320 294.800 ;
        RECT 19.730 268.200 71.790 284.200 ;
        RECT 10.870 262.800 71.790 268.200 ;
        RECT 10.870 260.200 54.370 262.800 ;
        RECT 2.800 252.200 54.370 260.200 ;
        RECT 2.800 246.800 72.200 252.200 ;
        RECT 2.800 230.800 57.850 246.800 ;
        RECT 4.120 228.200 57.850 230.800 ;
        RECT 4.120 214.800 71.790 228.200 ;
        RECT 11.615 206.800 71.790 214.800 ;
        RECT 11.615 204.200 64.565 206.800 ;
        RECT 2.800 198.800 64.565 204.200 ;
        RECT 10.840 196.200 64.565 198.800 ;
        RECT 10.840 134.800 71.790 196.200 ;
        RECT 10.840 132.200 70.155 134.800 ;
        RECT 4.785 124.200 70.155 132.200 ;
        RECT 4.110 118.800 70.635 124.200 ;
        RECT 4.110 116.200 59.035 118.800 ;
        RECT 2.800 68.200 59.035 116.200 ;
        RECT 1.000 46.800 74.000 68.200 ;
        RECT 1.000 18.200 23.200 46.800 ;
        RECT 51.800 18.200 74.000 46.800 ;
        RECT 1.000 0.000 74.000 18.200 ;
  END
END gf180mcu_fd_io__bi_24t
END LIBRARY

