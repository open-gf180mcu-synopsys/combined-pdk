magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< obsm1 >>
rect -32 13108 1032 69957
<< obsm2 >>
rect 0 49200 1000 65000
<< metal3 >>
rect 0 63600 230 65000
rect 782 63600 1000 65000
rect 0 49200 222 50600
rect 774 49200 1000 50600
<< obsm3 >>
rect 222 50960 782 63240
<< labels >>
rlabel metal3 s 774 49200 1000 50600 6 VSS
port 1 nsew ground bidirectional
rlabel metal3 s 782 63600 1000 65000 6 VSS
port 1 nsew ground bidirectional
rlabel metal3 s 0 63600 230 65000 6 VSS
port 1 nsew ground bidirectional
rlabel metal3 s 0 49200 222 50600 6 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string LEFclass PAD
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2932394
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2930508
<< end >>
