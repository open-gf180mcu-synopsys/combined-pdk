* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addf_1 A B CI S CO VDD VSS
X0 S a_161_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD CI a_195_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_195_21# B a_178_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_76_111# B a_59_21# VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD A a_76_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_178_21# A a_161_21# VSS nfet_03p3 w=0.85u l=0.3u
X6 a_59_21# CI a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X7 a_9_111# B VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 a_110_21# CI VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 VDD A a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X10 a_59_21# CI a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS B a_110_21# VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X13 CO a_59_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS CI a_195_21# VSS nfet_03p3 w=0.85u l=0.3u
X15 CO a_59_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 VSS A a_76_21# VSS nfet_03p3 w=0.85u l=0.3u
X17 a_161_21# a_59_21# a_110_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 a_76_21# B a_59_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 a_178_111# A a_161_21# VDD pfet_03p3 w=1.7u l=0.3u
X20 a_195_111# B a_178_111# VDD pfet_03p3 w=1.7u l=0.3u
X21 a_9_21# B VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 a_110_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X23 a_161_21# a_59_21# a_110_111# VDD pfet_03p3 w=1.7u l=0.3u
X24 a_110_111# CI VDD VDD pfet_03p3 w=1.7u l=0.3u
X25 VDD B a_110_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_110_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X27 S a_161_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addh_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addh_1 A B S CO VDD VSS
X0 VDD B a_19_16# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_19_16# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_19_16# CO VDD pfet_03p3 w=1.7u l=0.3u
X3 a_19_16# B a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 S a_91_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 VSS a_19_16# CO VSS nfet_03p3 w=0.85u l=0.3u
X6 S a_91_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_91_21# B a_91_111# VDD pfet_03p3 w=1.7u l=0.3u
X8 VDD a_19_16# a_91_21# VDD pfet_03p3 w=1.7u l=0.3u
X9 a_91_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 a_91_21# A a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 a_42_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_19_16# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X13 a_75_21# B a_91_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__and2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__and2_1 A B Y VDD VSS
X0 Y a_12_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD B a_12_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_12_21# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_12_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X4 a_28_21# A a_12_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 VSS B a_28_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__aoi21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__aoi21_1 A0 A1 B Y VDD VSS
X0 Y B a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_9_111# A1 VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD A0 a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS B Y VSS nfet_03p3 w=0.85u l=0.3u
X4 a_28_21# A0 VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A1 a_28_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__aoi22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__aoi22_1 Y A0 A1 B0 B1
X0 a_9_111# B1 Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y B0 a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_9_111# A1 VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD A0 a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X4 a_56_21# B0 Y VSS nfet_03p3 w=0.85u l=0.3u
X5 VSS B1 a_56_21# VSS nfet_03p3 w=0.85u l=0.3u
X6 a_28_21# A0 VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 Y A1 a_28_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_1 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_2 A Y VDD VSS
X0 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_4 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X6 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X8 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_8 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X6 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X8 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X9 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X10 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X11 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X15 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X17 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_16 A Y VDD VSS
X0 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X5 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X7 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X10 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X13 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X15 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X19 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X21 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X22 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X23 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X24 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X26 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X27 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X28 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X29 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X30 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X32 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X33 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
C0 VDD Y 2.003100fF
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_1 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_2 A Y VDD VSS
X0 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_4 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X6 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X8 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_8 A Y VDD VSS
X0 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X6 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X8 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X9 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X10 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X11 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X15 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X17 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_16 A Y VDD VSS
X0 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X3 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X5 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X7 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X10 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X13 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X15 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X19 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X21 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X22 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X23 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X24 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 Y a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X26 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X27 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X28 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X29 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X30 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 VDD a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X32 Y a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X33 VSS a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
C0 VDD Y 2.003150fF
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_1 A Y VDD VSS
X0 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_2 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_4 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_8 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X8 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X13 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X14 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X15 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_16 A Y VDD VSS
X0 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X6 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X8 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X9 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X16 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X19 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X20 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X21 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X22 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X23 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X24 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X25 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X26 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X27 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X28 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X29 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X31 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dff_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dff_1 D Q QN CLK VDD VSS
X0 a_19_16# CLK a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_75_111# a_52_16# a_19_16# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_135_70# a_114_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X4 a_131_21# a_52_16# a_114_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_42_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 a_135_70# a_114_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 VDD a_19_16# a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X8 a_75_21# CLK a_19_16# VSS nfet_03p3 w=0.85u l=0.3u
X9 VSS a_135_70# a_131_21# VSS nfet_03p3 w=0.85u l=0.3u
X10 a_19_16# a_52_16# a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_19_16# a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X12 a_52_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 VDD a_135_70# a_131_111# VDD pfet_03p3 w=1.7u l=0.3u
X14 a_131_111# CLK a_114_21# VDD pfet_03p3 w=1.7u l=0.3u
X15 VSS a_135_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X16 a_114_21# a_52_16# a_103_111# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_114_21# CLK a_103_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 a_52_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X19 a_42_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 VDD a_9_21# a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X21 a_103_111# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 a_103_21# a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X23 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X24 VSS a_9_21# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X25 VDD a_135_70# QN VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffn_1 Q QN D CLK VDD VSS
X0 a_19_16# a_52_83# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_75_111# a_52_16# a_19_16# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_131_21# a_52_16# a_114_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_42_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD a_19_16# a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X5 VDD a_135_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X6 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_75_21# a_52_83# a_19_16# VSS nfet_03p3 w=0.85u l=0.3u
X8 VSS a_135_70# a_131_21# VSS nfet_03p3 w=0.85u l=0.3u
X9 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_19_16# a_52_16# a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_19_16# a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_135_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X13 a_52_16# a_52_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X14 VDD a_135_70# a_131_111# VDD pfet_03p3 w=1.7u l=0.3u
X15 VSS CLK a_52_83# VSS nfet_03p3 w=0.85u l=0.3u
X16 a_131_111# a_52_83# a_114_21# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_114_21# a_52_16# a_103_111# VDD pfet_03p3 w=1.7u l=0.3u
X18 a_114_21# a_52_83# a_103_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 a_135_70# a_114_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X20 a_52_16# a_52_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
X21 a_42_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 VDD a_9_21# a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_103_111# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X24 a_103_21# a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 a_135_70# a_114_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X26 VSS a_9_21# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X27 VDD CLK a_52_83# VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffr_1 D Q QN CLK RN VDD VSS
X0 a_122_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_205_70# a_201_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_62_100# CLK a_112_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 a_145_111# a_122_16# a_62_100# VDD pfet_03p3 w=1.7u l=0.3u
X4 a_145_21# CLK a_62_100# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 a_62_100# a_122_16# a_112_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_112_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X9 a_205_70# a_184_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 VDD a_205_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X12 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 a_201_21# a_122_16# a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS a_205_70# a_201_21# VSS nfet_03p3 w=0.85u l=0.3u
X15 a_205_70# a_25_21# a_273_111# VDD pfet_03p3 w=1.7u l=0.3u
X16 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 VSS a_205_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X18 a_273_111# a_184_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X19 VDD a_62_100# a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X20 VSS a_62_100# a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_112_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_173_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X24 VSS a_25_21# a_205_70# VSS nfet_03p3 w=0.85u l=0.3u
X25 a_201_111# CLK a_184_21# VDD pfet_03p3 w=1.7u l=0.3u
X26 VSS a_41_111# a_145_21# VSS nfet_03p3 w=0.85u l=0.3u
X27 a_184_21# a_122_16# a_173_111# VDD pfet_03p3 w=1.7u l=0.3u
X28 a_184_21# CLK a_173_21# VSS nfet_03p3 w=0.85u l=0.3u
X29 VDD a_41_111# a_145_111# VDD pfet_03p3 w=1.7u l=0.3u
X30 a_173_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 a_122_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffrn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffrn_1 D Q QN RN CLK VDD VSS
X0 a_122_16# a_122_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_205_70# a_201_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_62_100# a_122_83# a_112_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 a_145_111# a_122_16# a_62_100# VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS a_205_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X5 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 VDD a_205_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X7 a_145_21# a_122_83# a_62_100# VSS nfet_03p3 w=0.85u l=0.3u
X8 VSS a_25_21# a_205_70# VSS nfet_03p3 w=0.85u l=0.3u
X9 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 VDD CLK a_122_83# VDD pfet_03p3 w=1.7u l=0.3u
X11 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 a_62_100# a_122_16# a_112_21# VSS nfet_03p3 w=0.85u l=0.3u
X13 VSS CLK a_122_83# VSS nfet_03p3 w=0.85u l=0.3u
X14 a_205_70# a_184_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X15 a_112_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 a_201_21# a_122_16# a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS a_205_70# a_201_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 a_205_70# a_25_21# a_306_111# VDD pfet_03p3 w=1.7u l=0.3u
X21 a_306_111# a_184_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 VDD a_62_100# a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 VSS a_62_100# a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X24 a_112_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_173_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X27 a_201_111# a_122_83# a_184_21# VDD pfet_03p3 w=1.7u l=0.3u
X28 VSS a_41_111# a_145_21# VSS nfet_03p3 w=0.85u l=0.3u
X29 a_184_21# a_122_16# a_173_111# VDD pfet_03p3 w=1.7u l=0.3u
X30 a_184_21# a_122_83# a_173_21# VSS nfet_03p3 w=0.85u l=0.3u
X31 VDD a_41_111# a_145_111# VDD pfet_03p3 w=1.7u l=0.3u
X32 a_173_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X33 a_122_16# a_122_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffs_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffs_1 D Q QN SN CLK VDD VSS
X0 a_75_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X2 VSS SN a_108_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_227_21# a_147_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X4 a_208_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 VDD a_147_21# a_208_111# VDD pfet_03p3 w=1.7u l=0.3u
X6 a_85_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 a_168_70# SN a_227_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_85_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X9 a_75_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VDD a_168_70# a_164_111# VDD pfet_03p3 w=1.7u l=0.3u
X11 VDD SN SN VDD pfet_03p3 w=1.7u l=0.3u
X12 SN a_34_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 a_147_21# a_85_16# a_136_111# VDD pfet_03p3 w=1.7u l=0.3u
X14 a_164_111# CLK a_147_21# VDD pfet_03p3 w=1.7u l=0.3u
X15 a_136_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 VDD SN a_108_111# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_136_21# SN VSS VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS a_168_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X19 a_164_21# a_85_16# a_147_21# VSS nfet_03p3 w=0.85u l=0.3u
X20 a_108_111# a_85_16# a_34_16# VDD pfet_03p3 w=1.7u l=0.3u
X21 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 a_147_21# CLK a_136_21# VSS nfet_03p3 w=0.85u l=0.3u
X23 VDD a_168_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X24 VSS a_168_70# a_164_21# VSS nfet_03p3 w=0.85u l=0.3u
X25 a_34_16# CLK a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_29_21# SN SN VSS nfet_03p3 w=0.85u l=0.3u
X27 a_34_16# a_85_16# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X28 VSS a_34_16# a_29_21# VSS nfet_03p3 w=0.85u l=0.3u
X29 a_108_21# CLK a_34_16# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsn_1 D Q QN CLK SN VDD VSS
X0 a_75_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_147_21# a_242_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_242_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS SN a_108_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS CLK a_85_83# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_85_16# a_85_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_85_16# a_85_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_75_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X8 VDD a_168_70# a_164_111# VDD pfet_03p3 w=1.7u l=0.3u
X9 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VDD SN SN VDD pfet_03p3 w=1.7u l=0.3u
X11 SN a_34_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X12 a_147_21# a_85_16# a_136_111# VDD pfet_03p3 w=1.7u l=0.3u
X13 a_164_111# a_85_83# a_147_21# VDD pfet_03p3 w=1.7u l=0.3u
X14 VDD CLK a_85_83# VDD pfet_03p3 w=1.7u l=0.3u
X15 a_261_21# a_147_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 VSS a_168_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X17 a_136_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X18 VDD SN a_108_111# VDD pfet_03p3 w=1.7u l=0.3u
X19 a_136_21# SN VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 a_164_21# a_85_16# a_147_21# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_168_70# SN a_261_21# VSS nfet_03p3 w=0.85u l=0.3u
X22 a_108_111# a_85_16# a_34_16# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_147_21# a_85_83# a_136_21# VSS nfet_03p3 w=0.85u l=0.3u
X24 VSS a_168_70# a_164_21# VSS nfet_03p3 w=0.85u l=0.3u
X25 a_34_16# a_85_83# a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_29_21# SN SN VSS nfet_03p3 w=0.85u l=0.3u
X27 a_34_16# a_85_16# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X28 VDD a_168_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X29 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 VSS a_34_16# a_29_21# VSS nfet_03p3 w=0.85u l=0.3u
X31 a_108_21# a_85_83# a_34_16# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsr_1 D Q QN RN SN CLK VDD VSS
X0 a_82_16# CLK a_123_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_212_111# CLK a_195_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS a_41_111# a_156_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_195_21# CLK a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS a_25_21# a_216_70# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_133_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_216_70# SN a_275_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 a_123_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 VDD a_216_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X9 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X11 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 a_82_16# a_133_16# a_123_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 a_256_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X15 a_275_21# a_195_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 VDD a_195_21# a_256_111# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_212_21# a_133_16# a_195_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 a_216_70# a_25_21# a_256_111# VDD pfet_03p3 w=1.7u l=0.3u
X19 VSS a_216_70# a_212_21# VSS nfet_03p3 w=0.85u l=0.3u
X20 a_77_21# SN a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_57_111# a_82_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 VDD SN a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X24 a_195_21# a_133_16# a_184_111# VDD pfet_03p3 w=1.7u l=0.3u
X25 VSS a_82_16# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X26 a_156_21# CLK a_82_16# VSS nfet_03p3 w=0.85u l=0.3u
X27 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X28 VDD a_41_111# a_156_111# VDD pfet_03p3 w=1.7u l=0.3u
X29 a_184_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 a_133_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 a_123_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X32 a_184_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X33 VSS a_216_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X34 a_156_111# a_133_16# a_82_16# VDD pfet_03p3 w=1.7u l=0.3u
X35 VDD a_216_70# a_212_111# VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsrn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsrn_1 D Q QN CLK RN SN VDD VSS
X0 a_82_16# a_133_83# a_123_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_212_111# a_133_83# a_195_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD CLK a_133_83# VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS a_41_111# a_156_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 a_195_21# a_133_83# a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_133_16# a_133_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_123_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 VSS a_216_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X10 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X11 a_310_21# a_195_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 VDD a_216_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X13 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 a_82_16# a_133_16# a_123_21# VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS CLK a_133_83# VSS nfet_03p3 w=0.85u l=0.3u
X16 a_216_70# SN a_310_21# VSS nfet_03p3 w=0.85u l=0.3u
X17 a_212_21# a_133_16# a_195_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS a_216_70# a_212_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 a_77_21# SN a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X20 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X21 a_57_111# a_82_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 a_216_70# a_25_21# a_291_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X24 VDD SN a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X25 a_195_21# a_133_16# a_184_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 VDD a_195_21# a_291_111# VDD pfet_03p3 w=1.7u l=0.3u
X27 a_291_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X28 VSS a_82_16# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X29 a_156_21# a_133_83# a_82_16# VSS nfet_03p3 w=0.85u l=0.3u
X30 VDD a_41_111# a_156_111# VDD pfet_03p3 w=1.7u l=0.3u
X31 a_184_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X32 a_133_16# a_133_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X33 a_123_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X34 a_184_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X35 VSS a_25_21# a_216_70# VSS nfet_03p3 w=0.85u l=0.3u
X36 a_156_111# a_133_16# a_82_16# VDD pfet_03p3 w=1.7u l=0.3u
X37 VDD a_216_70# a_212_111# VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dlat_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dlat_1 D Q CLK VDD VSS
X0 a_52_94# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 a_46_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X2 a_20_16# CLK a_46_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 VSS a_10_21# a_127_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 a_77_111# CLK a_20_16# VDD pfet_03p3 w=1.7u l=0.3u
X5 VDD a_10_21# a_77_111# VDD pfet_03p3 w=1.7u l=0.3u
X6 a_20_16# a_52_94# a_43_111# VDD pfet_03p3 w=1.7u l=0.3u
X7 VDD a_20_16# a_10_21# VDD pfet_03p3 w=1.7u l=0.3u
X8 a_43_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X9 Q a_127_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 VDD a_10_21# a_127_21# VDD pfet_03p3 w=1.7u l=0.3u
X11 a_77_21# a_52_94# a_20_16# VSS nfet_03p3 w=0.85u l=0.3u
X12 Q a_127_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 VSS a_10_21# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 a_52_94# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS a_20_16# a_10_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dlatn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dlatn_1 D Q CLK VDD VSS
X0 VDD CLK a_54_16# VDD pfet_03p3 w=1.7u l=0.3u
X1 Q a_161_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X2 a_52_94# a_54_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS CLK a_54_16# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS a_10_21# a_161_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_46_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_20_16# a_54_16# a_46_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 a_77_111# a_54_16# a_20_16# VDD pfet_03p3 w=1.7u l=0.3u
X8 VDD a_10_21# a_77_111# VDD pfet_03p3 w=1.7u l=0.3u
X9 a_20_16# a_52_94# a_43_111# VDD pfet_03p3 w=1.7u l=0.3u
X10 VDD a_20_16# a_10_21# VDD pfet_03p3 w=1.7u l=0.3u
X11 a_43_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X12 Q a_161_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 VDD a_10_21# a_161_21# VDD pfet_03p3 w=1.7u l=0.3u
X14 a_77_21# a_52_94# a_20_16# VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS a_10_21# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X16 a_52_94# a_54_16# VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 VSS a_20_16# a_10_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_1 VDD VSS
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_2 VDD VSS
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_4 VDD VSS
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_8 VDD VSS
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_16 VDD VSS
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_1 A Y VDD VSS
X0 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_2 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_4 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X3 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X7 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_8 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X8 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X13 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X14 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X15 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_16 A Y VDD VSS
X0 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X6 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X8 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X9 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X16 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X18 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X19 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X20 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X21 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X22 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X23 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X24 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X25 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X26 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X27 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X28 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X29 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X31 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__lshifdown.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__lshifdown A Y VDDH VDD VSS
X0 a_26_21# A VDDH VDDH pfet_03p3 w=1.7u l=0.3u
X1 Y a_26_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X2 Y a_26_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 a_26_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__lshifup.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__lshifup A Y VDDH VDD VSS
X0 a_26_21# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_67_21# VDDH VDDH pfet_03p3 w=1.7u l=0.3u
X2 VSS A a_67_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 Y a_67_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X4 VDDH a_78_84# a_67_21# VDDH pfet_03p3 w=1.7u l=0.3u
X5 a_78_84# a_67_21# VDDH VDDH pfet_03p3 w=1.7u l=0.3u
X6 a_26_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 a_78_84# a_26_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__mux2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__mux2_1 A B Y Sel VDD VSS
X0 B a_25_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y Sel A VDD pfet_03p3 w=1.7u l=0.3u
X2 a_25_21# Sel VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 Y a_25_21# A VSS nfet_03p3 w=0.85u l=0.3u
X4 a_25_21# Sel VSS VSS nfet_03p3 w=0.85u l=0.3u
X5 B Sel Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nand2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__nand2_1 A B Y VDD VSS
X0 VDD B Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 a_28_21# A Y VSS nfet_03p3 w=0.85u l=0.3u
X3 VSS B a_28_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__nor2_1 A B Y VDD VSS
X0 Y B a_25_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_25_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 VSS B Y VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai21_1 A0 A1 B Y VDD VSS
X0 Y B a_8_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 VSS A0 a_8_21# VSS nfet_03p3 w=0.85u l=0.3u
X2 a_27_111# A0 VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD B Y VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A1 a_27_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_8_21# A1 VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai22_1 A0 A1 B0 B1 Y VDD VSS
X0 a_8_21# B1 Y VSS nfet_03p3 w=0.85u l=0.3u
X1 Y B0 a_8_21# VSS nfet_03p3 w=0.85u l=0.3u
X2 VSS A0 a_8_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 VDD B1 a_56_111# VDD pfet_03p3 w=1.7u l=0.3u
X4 a_27_111# A0 VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 a_56_111# B0 Y VDD pfet_03p3 w=1.7u l=0.3u
X6 Y A1 a_27_111# VDD pfet_03p3 w=1.7u l=0.3u
X7 a_8_21# A1 VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai31_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai31_1 A0 A1 A2 B Y VDD VSS
X0 a_35_111# A0 VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 a_25_21# A2 VSS VSS nfet_03p3 w=0.85u l=0.3u
X2 a_25_21# A0 VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 Y B a_25_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 Y A2 a_46_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 VDD B Y VDD pfet_03p3 w=1.7u l=0.3u
X6 VSS A1 a_25_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 a_46_111# A1 a_35_111# VDD pfet_03p3 w=1.7u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__or2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__or2_1 A B Y VDD VSS
X0 VDD B a_25_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_25_111# A a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 Y a_9_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 a_9_111# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X4 Y a_9_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS B a_9_111# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tbuf_1 A Y EN VDD VSS
X0 Y EN a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 Y a_47_96# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_42_111# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_47_96# EN VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_47_96# EN VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_42_21# a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tieh.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tieh Y VDD VSS
X0 Y a_19_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 a_19_16# a_19_16# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tiel.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tiel Y VDD VSS
X0 a_19_16# a_19_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 Y a_19_16# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tinv_1 A Y EN VDD VSS
X0 Y EN a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 Y a_9_21# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_42_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD EN a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS EN a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_42_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__xnor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__xnor2_1 A B Y VDD VSS
X0 Y a_47_16# a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 a_47_16# B VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD B a_76_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 a_76_111# A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 Y a_47_16# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_42_111# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X7 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_76_21# a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X9 a_42_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_47_16# B VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS B a_76_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__xor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__xor2_1 A B Y VDD VSS
X0 Y B a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 a_47_96# B VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD B a_76_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 a_76_111# a_9_21# Y VDD pfet_03p3 w=1.7u l=0.3u
X4 Y a_47_96# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_42_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 VDD A a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X7 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_76_21# a_9_21# Y VSS nfet_03p3 w=0.85u l=0.3u
X9 a_42_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_47_96# B VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_47_96# a_76_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends


******* EOF

