magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 1620 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 850 210 910 380
rect 1020 210 1080 380
rect 1190 210 1250 380
rect 1360 210 1420 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 530 1110 590 1450
rect 850 1110 910 1450
rect 1020 1110 1080 1450
rect 1190 1110 1250 1450
rect 1360 1110 1420 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 530 380
rect 590 318 690 380
rect 590 272 622 318
rect 668 272 690 318
rect 590 210 690 272
rect 750 318 850 380
rect 750 272 772 318
rect 818 272 850 318
rect 750 210 850 272
rect 910 358 1020 380
rect 910 312 942 358
rect 988 312 1020 358
rect 910 210 1020 312
rect 1080 318 1190 380
rect 1080 272 1112 318
rect 1158 272 1190 318
rect 1080 210 1190 272
rect 1250 318 1360 380
rect 1250 272 1282 318
rect 1328 272 1360 318
rect 1250 210 1360 272
rect 1420 318 1520 380
rect 1420 272 1452 318
rect 1498 272 1520 318
rect 1420 210 1520 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1397 530 1450
rect 420 1163 452 1397
rect 498 1163 530 1397
rect 420 1110 530 1163
rect 590 1397 690 1450
rect 590 1163 622 1397
rect 668 1163 690 1397
rect 590 1110 690 1163
rect 750 1397 850 1450
rect 750 1163 772 1397
rect 818 1163 850 1397
rect 750 1110 850 1163
rect 910 1110 1020 1450
rect 1080 1397 1190 1450
rect 1080 1163 1112 1397
rect 1158 1163 1190 1397
rect 1080 1110 1190 1163
rect 1250 1397 1360 1450
rect 1250 1163 1282 1397
rect 1328 1163 1360 1397
rect 1250 1110 1360 1163
rect 1420 1397 1520 1450
rect 1420 1163 1452 1397
rect 1498 1163 1520 1397
rect 1420 1110 1520 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 622 272 668 318
rect 772 272 818 318
rect 942 312 988 358
rect 1112 272 1158 318
rect 1282 272 1328 318
rect 1452 272 1498 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 452 1163 498 1397
rect 622 1163 668 1397
rect 772 1163 818 1397
rect 1112 1163 1158 1397
rect 1282 1163 1328 1397
rect 1452 1163 1498 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 300 1588 450 1610
rect 300 1542 352 1588
rect 398 1542 450 1588
rect 300 1520 450 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1020 1588 1170 1610
rect 1020 1542 1072 1588
rect 1118 1542 1170 1588
rect 1020 1520 1170 1542
rect 1260 1588 1410 1610
rect 1260 1542 1312 1588
rect 1358 1542 1410 1588
rect 1260 1520 1410 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 352 1542 398 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1072 1542 1118 1588
rect 1312 1542 1358 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 530 1450 590 1500
rect 850 1450 910 1500
rect 1020 1450 1080 1500
rect 1190 1450 1250 1500
rect 1360 1450 1420 1500
rect 190 1060 250 1110
rect 190 1033 310 1060
rect 190 987 237 1033
rect 283 987 310 1033
rect 190 960 310 987
rect 190 380 250 960
rect 360 800 420 1110
rect 300 773 420 800
rect 300 727 327 773
rect 373 727 420 773
rect 300 700 420 727
rect 360 380 420 700
rect 530 670 590 1110
rect 850 800 910 1110
rect 780 773 910 800
rect 780 727 807 773
rect 853 727 910 773
rect 780 700 910 727
rect 470 643 590 670
rect 470 597 497 643
rect 543 597 590 643
rect 470 570 590 597
rect 530 380 590 570
rect 850 380 910 700
rect 1020 670 1080 1110
rect 1190 1060 1250 1110
rect 1190 1033 1310 1060
rect 1190 987 1237 1033
rect 1283 987 1310 1033
rect 1190 960 1310 987
rect 1020 643 1140 670
rect 1020 597 1067 643
rect 1113 597 1140 643
rect 1020 570 1140 597
rect 1020 380 1080 570
rect 1190 380 1250 960
rect 1360 800 1420 1110
rect 1300 773 1420 800
rect 1300 727 1327 773
rect 1373 727 1420 773
rect 1300 700 1420 727
rect 1360 380 1420 700
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 850 160 910 210
rect 1020 160 1080 210
rect 1190 160 1250 210
rect 1360 160 1420 210
<< polycontact >>
rect 237 987 283 1033
rect 327 727 373 773
rect 807 727 853 773
rect 497 597 543 643
rect 1237 987 1283 1033
rect 1067 597 1113 643
rect 1327 727 1373 773
<< metal1 >>
rect 0 1588 1620 1660
rect 0 1542 112 1588
rect 158 1542 352 1588
rect 398 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1072 1588
rect 1118 1542 1312 1588
rect 1358 1542 1620 1588
rect 0 1520 1620 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 520 160 1163
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 450 1397 500 1450
rect 450 1163 452 1397
rect 498 1163 500 1397
rect 450 1040 500 1163
rect 620 1397 670 1520
rect 620 1163 622 1397
rect 668 1163 670 1397
rect 620 1110 670 1163
rect 770 1397 820 1520
rect 770 1163 772 1397
rect 818 1163 820 1397
rect 770 1110 820 1163
rect 1110 1397 1160 1450
rect 1110 1163 1112 1397
rect 1158 1163 1160 1397
rect 210 1036 700 1040
rect 210 1033 624 1036
rect 210 987 237 1033
rect 283 987 624 1033
rect 210 984 624 987
rect 676 984 700 1036
rect 210 980 700 984
rect 300 776 400 780
rect 300 724 324 776
rect 376 724 400 776
rect 300 720 400 724
rect 470 646 570 650
rect 470 594 494 646
rect 546 594 570 646
rect 470 590 570 594
rect 80 516 180 520
rect 80 464 104 516
rect 156 464 180 516
rect 80 460 180 464
rect 110 318 160 460
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 620 318 670 980
rect 1110 780 1160 1163
rect 1280 1397 1330 1520
rect 1280 1163 1282 1397
rect 1328 1163 1330 1397
rect 1280 1110 1330 1163
rect 1450 1397 1500 1450
rect 1450 1163 1452 1397
rect 1498 1163 1500 1397
rect 1450 1050 1500 1163
rect 1450 1040 1520 1050
rect 1210 1036 1310 1040
rect 1210 984 1234 1036
rect 1286 984 1310 1036
rect 1210 980 1310 984
rect 1440 1036 1540 1040
rect 1440 984 1464 1036
rect 1516 984 1540 1036
rect 1440 980 1540 984
rect 1450 970 1520 980
rect 780 776 880 780
rect 780 724 804 776
rect 856 724 880 776
rect 1110 773 1400 780
rect 1110 770 1327 773
rect 780 720 880 724
rect 940 727 1327 770
rect 1373 727 1400 773
rect 940 720 1400 727
rect 620 272 622 318
rect 668 272 670 318
rect 620 210 670 272
rect 770 318 820 400
rect 770 272 772 318
rect 818 272 820 318
rect 940 358 990 720
rect 1040 646 1140 650
rect 1040 594 1064 646
rect 1116 594 1140 646
rect 1040 590 1140 594
rect 940 312 942 358
rect 988 312 990 358
rect 940 290 990 312
rect 1110 318 1160 400
rect 770 240 820 272
rect 1110 272 1112 318
rect 1158 272 1160 318
rect 1110 240 1160 272
rect 770 190 1160 240
rect 1280 318 1330 380
rect 1280 272 1282 318
rect 1328 272 1330 318
rect 1280 140 1330 272
rect 1450 318 1500 970
rect 1450 272 1452 318
rect 1498 272 1500 318
rect 1450 210 1500 272
rect 0 118 1620 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1620 118
rect 0 0 1620 72
<< via1 >>
rect 624 984 676 1036
rect 324 773 376 776
rect 324 727 327 773
rect 327 727 373 773
rect 373 727 376 773
rect 324 724 376 727
rect 494 643 546 646
rect 494 597 497 643
rect 497 597 543 643
rect 543 597 546 643
rect 494 594 546 597
rect 104 464 156 516
rect 1234 1033 1286 1036
rect 1234 987 1237 1033
rect 1237 987 1283 1033
rect 1283 987 1286 1033
rect 1234 984 1286 987
rect 1464 984 1516 1036
rect 804 773 856 776
rect 804 727 807 773
rect 807 727 853 773
rect 853 727 856 773
rect 804 724 856 727
rect 1064 643 1116 646
rect 1064 597 1067 643
rect 1067 597 1113 643
rect 1113 597 1116 643
rect 1064 594 1116 597
<< metal2 >>
rect 600 1040 700 1050
rect 1210 1040 1310 1050
rect 600 1036 1310 1040
rect 600 984 624 1036
rect 676 984 1234 1036
rect 1286 984 1310 1036
rect 600 980 1310 984
rect 600 970 700 980
rect 1210 970 1310 980
rect 1440 1036 1540 1050
rect 1440 984 1464 1036
rect 1516 984 1540 1036
rect 1440 970 1540 984
rect 300 780 400 790
rect 780 780 880 790
rect 300 776 880 780
rect 300 724 324 776
rect 376 724 804 776
rect 856 724 880 776
rect 300 720 880 724
rect 300 710 400 720
rect 780 710 880 720
rect 470 650 570 660
rect 1040 650 1140 660
rect 470 646 1140 650
rect 470 594 494 646
rect 546 594 1064 646
rect 1116 594 1140 646
rect 470 590 1140 594
rect 470 580 570 590
rect 1040 580 1140 590
rect 80 516 180 530
rect 80 464 104 516
rect 156 464 180 516
rect 80 450 180 464
<< labels >>
rlabel via1 s 804 724 856 776 4 A
port 1 nsew signal input
rlabel via1 s 1064 594 1116 646 4 B
port 2 nsew signal input
rlabel via1 s 1464 984 1516 1036 4 S
port 3 nsew signal output
rlabel via1 s 104 464 156 516 4 CO
port 4 nsew signal output
rlabel metal1 s 280 1110 330 1660 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 620 1110 670 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 770 1110 820 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1280 1110 1330 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 1520 1620 1660 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1280 0 1330 380 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1620 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel via1 s 324 724 376 776 1 A
port 1 nsew signal input
rlabel metal2 s 300 710 400 790 1 A
port 1 nsew signal input
rlabel metal2 s 300 720 880 780 1 A
port 1 nsew signal input
rlabel metal2 s 780 710 880 790 1 A
port 1 nsew signal input
rlabel metal1 s 300 720 400 780 1 A
port 1 nsew signal input
rlabel metal1 s 780 720 880 780 1 A
port 1 nsew signal input
rlabel via1 s 494 594 546 646 1 B
port 2 nsew signal input
rlabel metal2 s 470 580 570 660 1 B
port 2 nsew signal input
rlabel metal2 s 470 590 1140 650 1 B
port 2 nsew signal input
rlabel metal2 s 1040 580 1140 660 1 B
port 2 nsew signal input
rlabel metal1 s 470 590 570 650 1 B
port 2 nsew signal input
rlabel metal1 s 1040 590 1140 650 1 B
port 2 nsew signal input
rlabel metal2 s 80 450 180 530 1 CO
port 4 nsew signal output
rlabel metal1 s 110 210 160 1450 1 CO
port 4 nsew signal output
rlabel metal1 s 80 460 180 520 1 CO
port 4 nsew signal output
rlabel metal2 s 1440 970 1540 1050 1 S
port 3 nsew signal output
rlabel metal1 s 1450 210 1500 1450 1 S
port 3 nsew signal output
rlabel metal1 s 1450 970 1520 1050 1 S
port 3 nsew signal output
rlabel metal1 s 1440 980 1540 1040 1 S
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1620 1660
string GDS_END 30160
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 19236
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
