magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use M1_NWELL05_512x8m81  M1_NWELL05_512x8m81_0
timestamp 1750858719
transform 1 0 310 0 1 12142
box 0 0 1 1
use M1_NWELL09_512x8m81  M1_NWELL09_512x8m81_0
timestamp 1750858719
transform 1 0 237 0 1 1392
box 0 0 1 1
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1750858719
transform 1 0 287 0 1 10310
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1750858719
transform 1 0 310 0 1 3446
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1750858719
transform 1 0 310 0 1 3169
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1750858719
transform 1 0 253 0 1 1202
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1750858719
transform 1 0 316 0 1 7141
box 0 0 1 1
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1750858719
transform 1 0 0 0 1 5237
box 0 0 1 1
use M1_PSUB$$47122476_512x8m81  M1_PSUB$$47122476_512x8m81_0
timestamp 1750858719
transform 1 0 237 0 1 73
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1750858719
transform 1 0 311 0 1 10780
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1750858719
transform 1 0 311 0 1 11555
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1750858719
transform 1 0 96 0 1 9560
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_3
timestamp 1750858719
transform 1 0 108 0 1 8520
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_4
timestamp 1750858719
transform 1 0 252 0 1 986
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_5
timestamp 1750858719
transform 1 0 316 0 1 7088
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_6
timestamp 1750858719
transform 1 0 526 0 1 9560
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1750858719
transform 1 0 394 0 1 5241
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1750858719
transform 1 0 101 0 1 5439
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_2
timestamp 1750858719
transform 1 0 312 0 1 1201
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_3
timestamp 1750858719
transform 1 0 310 0 1 3169
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_4
timestamp 1750858719
transform 1 0 526 0 1 5033
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_0
timestamp 1750858719
transform 1 0 394 0 1 5176
box 0 0 1 1
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_0
timestamp 1750858719
transform 1 0 281 0 -1 4915
box -31 0 -30 1
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_1
timestamp 1750858719
transform 1 0 281 0 -1 6919
box -31 0 -30 1
use nmos_5p0431059130202_512x8m81  nmos_5p0431059130202_512x8m81_0
timestamp 1750858719
transform 1 0 52 0 1 383
box 0 0 1 1
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_0
timestamp 1750858719
transform 1 0 281 0 -1 3060
box -31 0 -30 1
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1750858719
transform 1 0 248 0 -1 10197
box 0 0 1 1
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_1
timestamp 1750858719
transform 1 0 250 0 -1 8610
box 0 0 1 1
use via1_2_512x8m81  via1_2_512x8m81_0
timestamp 1750858719
transform 1 0 264 0 1 88
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1750858719
transform 0 -1 378 1 0 3387
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_1
timestamp 1750858719
transform 0 -1 373 1 0 12131
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1750858719
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1750858719
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_512x8m81  via2_R90_512x8m81_1
timestamp 1750858719
transform 0 -1 373 1 0 12131
box 0 0 1 1
<< properties >>
string GDS_END 307026
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 297780
string path 0.000 27.385 0.000 -0.005 
<< end >>
