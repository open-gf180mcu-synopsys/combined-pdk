magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1340 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 520 210 580 380
rect 750 210 810 380
rect 910 210 970 380
rect 1080 210 1140 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 520 720 580 1060
rect 750 720 810 1060
rect 910 720 970 1060
rect 1080 720 1140 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 520 380
rect 580 278 750 380
rect 580 232 642 278
rect 688 232 750 278
rect 580 210 750 232
rect 810 210 910 380
rect 970 313 1080 380
rect 970 267 1002 313
rect 1048 267 1080 313
rect 970 210 1080 267
rect 1140 318 1240 380
rect 1140 272 1172 318
rect 1218 272 1240 318
rect 1140 210 1240 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1037 360 1060
rect 250 803 282 1037
rect 328 803 360 1037
rect 250 720 360 803
rect 420 720 520 1060
rect 580 1038 750 1060
rect 580 992 642 1038
rect 688 992 750 1038
rect 580 720 750 992
rect 810 720 910 1060
rect 970 1037 1080 1060
rect 970 803 1002 1037
rect 1048 803 1080 1037
rect 970 720 1080 803
rect 1140 1007 1240 1060
rect 1140 773 1172 1007
rect 1218 773 1240 1007
rect 1140 720 1240 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 642 232 688 278
rect 1002 267 1048 313
rect 1172 272 1218 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 803 328 1037
rect 642 992 688 1038
rect 1002 803 1048 1037
rect 1172 773 1218 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 520 1060 580 1110
rect 750 1060 810 1110
rect 910 1060 970 1110
rect 1080 1060 1140 1110
rect 190 700 250 720
rect 360 700 420 720
rect 190 650 420 700
rect 520 700 580 720
rect 750 700 810 720
rect 520 678 620 700
rect 190 540 250 650
rect 520 632 547 678
rect 593 632 620 678
rect 520 610 620 632
rect 710 673 810 700
rect 710 627 737 673
rect 783 627 810 673
rect 910 700 970 720
rect 1080 700 1140 720
rect 910 650 1140 700
rect 710 600 810 627
rect 190 513 320 540
rect 190 467 247 513
rect 293 467 320 513
rect 190 440 320 467
rect 470 473 580 500
rect 190 400 420 440
rect 470 427 497 473
rect 543 427 580 473
rect 470 400 580 427
rect 190 380 250 400
rect 360 380 420 400
rect 520 380 580 400
rect 750 380 810 600
rect 870 578 970 600
rect 870 532 897 578
rect 943 532 970 578
rect 1080 540 1140 650
rect 870 510 970 532
rect 910 380 970 510
rect 1020 513 1140 540
rect 1020 467 1047 513
rect 1093 467 1140 513
rect 1020 440 1140 467
rect 1080 380 1140 440
rect 190 160 250 210
rect 360 160 420 210
rect 520 160 580 210
rect 750 160 810 210
rect 910 160 970 210
rect 1080 160 1140 210
<< polycontact >>
rect 547 632 593 678
rect 737 627 783 673
rect 247 467 293 513
rect 497 427 543 473
rect 897 532 943 578
rect 1047 467 1093 513
<< metal1 >>
rect 0 1198 1340 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1340 1198
rect 0 1130 1340 1152
rect 110 1007 160 1060
rect 110 773 112 1007
rect 158 773 160 1007
rect 280 1037 330 1130
rect 280 803 282 1037
rect 328 803 330 1037
rect 640 1038 690 1060
rect 640 992 642 1038
rect 688 992 690 1038
rect 640 930 690 992
rect 630 910 690 930
rect 1000 1037 1050 1130
rect 610 906 710 910
rect 610 854 634 906
rect 686 854 710 906
rect 610 850 710 854
rect 280 780 330 803
rect 1000 803 1002 1037
rect 1048 803 1050 1037
rect 110 670 160 773
rect 540 750 940 800
rect 1000 780 1050 803
rect 1170 1007 1220 1060
rect 540 680 600 750
rect 890 700 940 750
rect 1170 773 1172 1007
rect 1218 773 1220 1007
rect 1170 700 1220 773
rect 520 678 620 680
rect 110 620 470 670
rect 520 632 547 678
rect 593 632 620 678
rect 520 630 620 632
rect 730 673 790 700
rect 110 318 160 620
rect 410 580 470 620
rect 730 627 737 673
rect 783 627 790 673
rect 730 580 790 627
rect 890 640 1220 700
rect 890 590 950 640
rect 410 530 790 580
rect 870 578 970 590
rect 870 532 897 578
rect 943 532 970 578
rect 870 530 970 532
rect 220 516 320 520
rect 220 464 244 516
rect 296 464 320 516
rect 1020 516 1120 520
rect 1020 480 1044 516
rect 220 460 320 464
rect 470 473 1044 480
rect 470 427 497 473
rect 543 464 1044 473
rect 1096 464 1120 516
rect 543 460 1120 464
rect 543 427 1090 460
rect 470 420 1090 427
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 630 360 690 370
rect 280 272 282 318
rect 328 272 330 318
rect 610 356 710 360
rect 610 304 634 356
rect 686 304 710 356
rect 610 300 710 304
rect 1000 313 1050 370
rect 630 280 690 300
rect 280 140 330 272
rect 640 278 690 280
rect 640 232 642 278
rect 688 232 690 278
rect 640 210 690 232
rect 1000 267 1002 313
rect 1048 267 1050 313
rect 1000 140 1050 267
rect 1170 318 1220 640
rect 1170 272 1172 318
rect 1218 272 1220 318
rect 1170 210 1220 272
rect 0 118 1340 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1340 118
rect 0 0 1340 72
<< via1 >>
rect 634 854 686 906
rect 244 513 296 516
rect 244 467 247 513
rect 247 467 293 513
rect 293 467 296 513
rect 244 464 296 467
rect 1044 513 1096 516
rect 1044 467 1047 513
rect 1047 467 1093 513
rect 1093 467 1096 513
rect 1044 464 1096 467
rect 634 304 686 356
<< metal2 >>
rect 630 920 690 930
rect 620 906 700 920
rect 620 854 634 906
rect 686 854 700 906
rect 620 840 700 854
rect 230 520 310 530
rect 220 516 320 520
rect 220 464 244 516
rect 296 464 320 516
rect 220 460 320 464
rect 230 450 310 460
rect 630 370 690 840
rect 1030 520 1110 530
rect 1020 516 1120 520
rect 1020 464 1044 516
rect 1096 464 1120 516
rect 1020 460 1120 464
rect 1030 450 1110 460
rect 610 356 710 370
rect 610 304 634 356
rect 686 304 710 356
rect 610 290 710 304
<< labels >>
rlabel via1 s 244 464 296 516 4 A
port 1 nsew signal input
rlabel via1 s 1044 464 1096 516 4 B
port 2 nsew signal input
rlabel via1 s 634 304 686 356 4 Y
port 3 nsew signal output
rlabel metal1 s 280 780 330 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1000 780 1050 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1340 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1000 0 1050 370 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1340 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 230 450 310 530 1 A
port 1 nsew signal input
rlabel metal2 s 220 460 320 520 1 A
port 1 nsew signal input
rlabel metal1 s 220 460 320 520 1 A
port 1 nsew signal input
rlabel metal2 s 1030 450 1110 530 1 B
port 2 nsew signal input
rlabel metal2 s 1020 460 1120 520 1 B
port 2 nsew signal input
rlabel metal1 s 470 420 1090 480 1 B
port 2 nsew signal input
rlabel metal1 s 1020 460 1120 520 1 B
port 2 nsew signal input
rlabel via1 s 634 854 686 906 1 Y
port 3 nsew signal output
rlabel metal2 s 630 290 690 930 1 Y
port 3 nsew signal output
rlabel metal2 s 620 840 700 920 1 Y
port 3 nsew signal output
rlabel metal2 s 610 290 710 370 1 Y
port 3 nsew signal output
rlabel metal1 s 630 850 690 930 1 Y
port 3 nsew signal output
rlabel metal1 s 640 850 690 1060 1 Y
port 3 nsew signal output
rlabel metal1 s 610 850 710 910 1 Y
port 3 nsew signal output
rlabel metal1 s 640 210 690 370 1 Y
port 3 nsew signal output
rlabel metal1 s 630 280 690 370 1 Y
port 3 nsew signal output
rlabel metal1 s 610 300 710 360 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1340 1270
string GDS_END 395898
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 387252
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
