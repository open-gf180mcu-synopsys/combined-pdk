VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__bi_t
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_fd_io__bi_t ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 264.460 69.780 350.000 ;
    END
  END A
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 328.545 3.740 350.000 ;
    END
  END CS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 72.600 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 49.445 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 67.195 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.590 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 4.575 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 17.930 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 9.070 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 17.930 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 17.930 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 9.815 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 2.320 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 8.810 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 8.905 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 8.905 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 8.810 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 2.230 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 62.215 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 71.890 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 66.125 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 59.650 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 55.255 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 54.080 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 63.600 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 68.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 9.320 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 9.320 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 25.555 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 22.880 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 2.965 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
  END DVSS
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.385 334.920 11.765 350.000 ;
    END
  END IE
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 7.776000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 266.340 70.510 350.000 ;
    END
  END OE
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 258.720001 ;
    PORT
      LAYER Metal3 ;
        RECT 25.000 20.000 50.000 45.000 ;
    END
  END PAD
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.330 330.100 10.710 350.000 ;
    END
  END PD
  PIN PDRV0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.110 264.665 7.490 350.000 ;
    END
  END PDRV0
  PIN PDRV1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.820 264.990 8.200 350.000 ;
    END
  END PDRV1
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.350000 ;
    ANTENNADIFFAREA 2.980000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.965 330.420 6.345 350.000 ;
    END
  END PU
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.670 265.140 69.050 350.000 ;
    END
  END SL
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 56.170 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 71.290 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.800000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.860 319.900 71.240 350.000 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 328.245 3.060 348.375 ;
        RECT 4.040 330.120 5.665 348.375 ;
        RECT 6.645 330.120 6.810 348.375 ;
        RECT 4.040 328.245 6.810 330.120 ;
        RECT 0.000 264.365 6.810 328.245 ;
        RECT 8.500 329.800 10.030 348.375 ;
        RECT 11.010 334.620 11.085 348.375 ;
        RECT 12.065 334.620 68.370 348.375 ;
        RECT 11.010 329.800 68.370 334.620 ;
        RECT 8.500 264.840 68.370 329.800 ;
        RECT 71.540 319.600 75.000 348.375 ;
        RECT 70.810 266.040 75.000 319.600 ;
        RECT 8.500 264.690 69.100 264.840 ;
        RECT 7.790 264.365 69.100 264.690 ;
        RECT 0.000 264.160 69.100 264.365 ;
        RECT 70.080 264.160 75.000 266.040 ;
        RECT 0.000 0.000 75.000 264.160 ;
      LAYER Metal3 ;
        RECT 11.120 340.200 66.200 348.390 ;
        RECT 6.375 334.800 71.790 340.200 ;
        RECT 11.120 324.200 61.800 334.800 ;
        RECT 2.800 318.800 72.200 324.200 ;
        RECT 2.800 310.800 69.490 318.800 ;
        RECT 27.355 300.200 52.280 310.800 ;
        RECT 19.730 294.800 71.790 300.200 ;
        RECT 24.680 286.800 53.455 294.800 ;
        RECT 24.680 284.200 47.645 286.800 ;
        RECT 19.730 276.200 47.645 284.200 ;
        RECT 19.730 268.200 65.395 276.200 ;
        RECT 10.870 262.800 71.790 268.200 ;
        RECT 10.870 260.200 54.370 262.800 ;
        RECT 2.800 252.200 54.370 260.200 ;
        RECT 2.800 246.800 72.200 252.200 ;
        RECT 2.800 230.800 57.850 246.800 ;
        RECT 4.120 228.200 57.850 230.800 ;
        RECT 4.120 214.800 71.790 228.200 ;
        RECT 11.615 206.800 71.790 214.800 ;
        RECT 11.615 204.200 64.325 206.800 ;
        RECT 2.800 198.800 64.325 204.200 ;
        RECT 10.610 196.200 64.325 198.800 ;
        RECT 10.610 182.800 71.790 196.200 ;
        RECT 10.705 148.200 71.790 182.800 ;
        RECT 10.610 134.800 71.790 148.200 ;
        RECT 10.610 132.200 70.090 134.800 ;
        RECT 4.765 124.200 70.090 132.200 ;
        RECT 4.030 118.800 70.800 124.200 ;
        RECT 4.030 116.200 60.415 118.800 ;
        RECT 2.800 68.200 60.415 116.200 ;
        RECT 0.665 46.800 74.000 68.200 ;
        RECT 0.665 18.200 23.200 46.800 ;
        RECT 51.800 18.200 74.000 46.800 ;
        RECT 0.665 0.000 74.000 18.200 ;
  END
END gf180mcu_fd_io__bi_t
END LIBRARY

