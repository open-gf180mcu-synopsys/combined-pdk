magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 377 3782 870
rect -86 352 2122 377
rect 2342 352 3782 377
<< pwell >>
rect 2122 352 2342 377
rect -86 -86 3782 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 572 93 692 165
rect 796 93 916 165
rect 980 93 1100 165
rect 1348 93 1468 165
rect 1532 93 1652 165
rect 1792 68 1912 232
rect 2016 68 2136 232
rect 2328 68 2448 232
rect 2696 68 2816 232
rect 2920 68 3040 232
rect 3144 68 3264 232
rect 3368 68 3488 232
<< mvpmos >>
rect 144 524 244 596
rect 348 524 448 596
rect 592 519 692 596
rect 796 519 896 596
rect 1000 519 1100 596
rect 1348 497 1448 569
rect 1552 497 1652 569
rect 1812 497 1912 716
rect 2026 497 2126 716
rect 2328 497 2428 716
rect 2716 472 2816 716
rect 2930 472 3030 716
rect 3154 472 3254 716
rect 3368 472 3468 716
<< mvndiff >>
rect 2196 244 2268 257
rect 2196 232 2209 244
rect 1712 165 1792 232
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 572 165
rect 468 106 497 152
rect 543 106 572 152
rect 468 93 572 106
rect 692 152 796 165
rect 692 106 721 152
rect 767 106 796 152
rect 692 93 796 106
rect 916 93 980 165
rect 1100 152 1188 165
rect 1100 106 1129 152
rect 1175 106 1188 152
rect 1100 93 1188 106
rect 1260 152 1348 165
rect 1260 106 1273 152
rect 1319 106 1348 152
rect 1260 93 1348 106
rect 1468 93 1532 165
rect 1652 152 1792 165
rect 1652 106 1681 152
rect 1727 106 1792 152
rect 1652 93 1792 106
rect 1712 68 1792 93
rect 1912 152 2016 232
rect 1912 106 1941 152
rect 1987 106 2016 152
rect 1912 68 2016 106
rect 2136 198 2209 232
rect 2255 232 2268 244
rect 2255 198 2328 232
rect 2136 68 2328 198
rect 2448 152 2536 232
rect 2448 106 2477 152
rect 2523 106 2536 152
rect 2448 68 2536 106
rect 2608 192 2696 232
rect 2608 146 2621 192
rect 2667 146 2696 192
rect 2608 68 2696 146
rect 2816 152 2920 232
rect 2816 106 2845 152
rect 2891 106 2920 152
rect 2816 68 2920 106
rect 3040 192 3144 232
rect 3040 146 3069 192
rect 3115 146 3144 192
rect 3040 68 3144 146
rect 3264 155 3368 232
rect 3264 109 3293 155
rect 3339 109 3368 155
rect 3264 68 3368 109
rect 3488 191 3576 232
rect 3488 145 3517 191
rect 3563 145 3576 191
rect 3488 68 3576 145
<< mvpdiff >>
rect 1712 703 1812 716
rect 56 583 144 596
rect 56 537 69 583
rect 115 537 144 583
rect 56 524 144 537
rect 244 524 348 596
rect 448 583 592 596
rect 448 537 477 583
rect 523 537 592 583
rect 448 524 592 537
rect 512 519 592 524
rect 692 583 796 596
rect 692 537 721 583
rect 767 537 796 583
rect 692 519 796 537
rect 896 583 1000 596
rect 896 537 925 583
rect 971 537 1000 583
rect 896 519 1000 537
rect 1100 582 1188 596
rect 1100 536 1129 582
rect 1175 536 1188 582
rect 1712 569 1725 703
rect 1100 519 1188 536
rect 1260 556 1348 569
rect 1260 510 1273 556
rect 1319 510 1348 556
rect 1260 497 1348 510
rect 1448 556 1552 569
rect 1448 510 1477 556
rect 1523 510 1552 556
rect 1448 497 1552 510
rect 1652 563 1725 569
rect 1771 563 1812 703
rect 1652 497 1812 563
rect 1912 609 2026 716
rect 1912 563 1951 609
rect 1997 563 2026 609
rect 1912 497 2026 563
rect 2126 497 2328 716
rect 2428 703 2516 716
rect 2428 657 2457 703
rect 2503 657 2516 703
rect 2428 497 2516 657
rect 2628 639 2716 716
rect 2628 499 2641 639
rect 2687 499 2716 639
rect 2628 472 2716 499
rect 2816 661 2930 716
rect 2816 615 2845 661
rect 2891 615 2930 661
rect 2816 472 2930 615
rect 3030 639 3154 716
rect 3030 499 3079 639
rect 3125 499 3154 639
rect 3030 472 3154 499
rect 3254 661 3368 716
rect 3254 615 3283 661
rect 3329 615 3368 661
rect 3254 472 3368 615
rect 3468 639 3556 716
rect 3468 499 3497 639
rect 3543 499 3556 639
rect 3468 472 3556 499
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 497 106 543 152
rect 721 106 767 152
rect 1129 106 1175 152
rect 1273 106 1319 152
rect 1681 106 1727 152
rect 1941 106 1987 152
rect 2209 198 2255 244
rect 2477 106 2523 152
rect 2621 146 2667 192
rect 2845 106 2891 152
rect 3069 146 3115 192
rect 3293 109 3339 155
rect 3517 145 3563 191
<< mvpdiffc >>
rect 69 537 115 583
rect 477 537 523 583
rect 721 537 767 583
rect 925 537 971 583
rect 1129 536 1175 582
rect 1273 510 1319 556
rect 1477 510 1523 556
rect 1725 563 1771 703
rect 1951 563 1997 609
rect 2457 657 2503 703
rect 2641 499 2687 639
rect 2845 615 2891 661
rect 3079 499 3125 639
rect 3283 615 3329 661
rect 3497 499 3543 639
<< polysilicon >>
rect 1812 716 1912 760
rect 2026 716 2126 760
rect 2328 716 2428 760
rect 2716 716 2816 760
rect 2930 716 3030 760
rect 3154 716 3254 760
rect 3368 716 3468 760
rect 144 596 244 640
rect 348 596 448 640
rect 592 596 692 640
rect 796 596 896 640
rect 1000 596 1100 640
rect 144 477 244 524
rect 144 337 174 477
rect 220 337 244 477
rect 144 209 244 337
rect 124 165 244 209
rect 348 304 448 524
rect 1348 569 1448 613
rect 1552 569 1652 613
rect 348 258 387 304
rect 433 258 448 304
rect 348 209 448 258
rect 592 399 692 519
rect 592 353 617 399
rect 663 353 692 399
rect 592 209 692 353
rect 348 165 468 209
rect 572 165 692 209
rect 796 304 896 519
rect 796 258 815 304
rect 861 258 896 304
rect 796 209 896 258
rect 1000 358 1100 519
rect 1000 312 1013 358
rect 1059 312 1100 358
rect 1000 209 1100 312
rect 796 165 916 209
rect 980 165 1100 209
rect 1348 427 1448 497
rect 1348 287 1377 427
rect 1423 287 1448 427
rect 1348 209 1448 287
rect 1552 417 1652 497
rect 1552 371 1593 417
rect 1639 371 1652 417
rect 1552 209 1652 371
rect 1812 316 1912 497
rect 1812 276 1836 316
rect 1792 270 1836 276
rect 1882 270 1912 316
rect 2026 417 2126 497
rect 2026 371 2050 417
rect 2096 371 2126 417
rect 2026 276 2126 371
rect 2328 420 2428 497
rect 2328 374 2353 420
rect 2399 374 2428 420
rect 2328 276 2428 374
rect 2716 413 2816 472
rect 2716 367 2740 413
rect 2786 367 2816 413
rect 2716 357 2816 367
rect 2930 413 3030 472
rect 2930 367 2959 413
rect 3005 367 3030 413
rect 2930 357 3030 367
rect 3154 413 3254 472
rect 3154 367 3182 413
rect 3228 367 3254 413
rect 3154 357 3254 367
rect 3368 413 3468 472
rect 3368 367 3387 413
rect 3433 367 3468 413
rect 3368 357 3468 367
rect 2716 311 3468 357
rect 2716 276 2816 311
rect 1792 232 1912 270
rect 2016 232 2136 276
rect 1348 165 1468 209
rect 1532 165 1652 209
rect 124 49 244 93
rect 348 49 468 93
rect 572 49 692 93
rect 796 49 916 93
rect 980 49 1100 93
rect 1348 49 1468 93
rect 1532 49 1652 93
rect 2328 232 2448 276
rect 2696 232 2816 276
rect 2920 232 3040 311
rect 3144 232 3264 311
rect 3368 276 3468 311
rect 3368 232 3488 276
rect 1792 24 1912 68
rect 2016 24 2136 68
rect 2328 24 2448 68
rect 2696 24 2816 68
rect 2920 24 3040 68
rect 3144 24 3264 68
rect 3368 24 3488 68
<< polycontact >>
rect 174 337 220 477
rect 387 258 433 304
rect 617 353 663 399
rect 815 258 861 304
rect 1013 312 1059 358
rect 1377 287 1423 427
rect 1593 371 1639 417
rect 1836 270 1882 316
rect 2050 371 2096 417
rect 2353 374 2399 420
rect 2740 367 2786 413
rect 2959 367 3005 413
rect 3182 367 3228 413
rect 3387 367 3433 413
<< metal1 >>
rect 0 724 3696 844
rect 69 583 115 596
rect 466 583 534 724
rect 69 271 115 537
rect 173 491 420 542
rect 466 537 477 583
rect 523 537 534 583
rect 710 632 1175 678
rect 710 583 778 632
rect 710 537 721 583
rect 767 537 778 583
rect 914 537 925 583
rect 971 537 1074 583
rect 173 477 775 491
rect 173 337 174 477
rect 220 445 775 477
rect 220 337 221 445
rect 729 419 775 445
rect 1028 452 1074 537
rect 1129 582 1175 632
rect 1129 522 1175 536
rect 1273 556 1319 724
rect 1714 703 1782 724
rect 1273 497 1319 510
rect 1377 628 1641 678
rect 173 320 221 337
rect 270 353 617 399
rect 663 353 682 399
rect 729 364 979 419
rect 1028 405 1187 452
rect 923 358 979 364
rect 270 271 316 353
rect 923 312 1013 358
rect 1059 312 1072 358
rect 69 224 316 271
rect 376 304 872 307
rect 376 258 387 304
rect 433 258 815 304
rect 861 258 872 304
rect 1141 261 1187 405
rect 1377 427 1423 628
rect 1377 261 1423 287
rect 376 253 872 258
rect 167 152 217 224
rect 1007 215 1423 261
rect 1477 556 1523 569
rect 1477 317 1523 510
rect 1594 515 1641 628
rect 1714 563 1725 703
rect 1771 563 1782 703
rect 2446 703 2514 724
rect 2446 657 2457 703
rect 2503 657 2514 703
rect 2605 639 2701 663
rect 1927 609 2515 610
rect 1927 563 1951 609
rect 1997 563 2515 609
rect 1714 561 1782 563
rect 1594 469 2399 515
rect 1582 417 2120 423
rect 1582 371 1593 417
rect 1639 371 2050 417
rect 2096 371 2120 417
rect 1582 364 2120 371
rect 2353 420 2399 469
rect 2353 339 2399 374
rect 2469 419 2515 563
rect 2605 499 2641 639
rect 2687 536 2701 639
rect 2845 661 2891 724
rect 2845 588 2891 615
rect 3053 639 3138 663
rect 3053 536 3079 639
rect 2687 499 3079 536
rect 3125 536 3138 639
rect 3283 661 3329 724
rect 3283 588 3329 615
rect 3474 639 3563 665
rect 3474 536 3497 639
rect 3125 499 3497 536
rect 3543 499 3563 639
rect 2605 472 3563 499
rect 2469 413 3445 419
rect 2469 367 2740 413
rect 2786 367 2959 413
rect 3005 367 3182 413
rect 3228 367 3387 413
rect 3433 367 3445 413
rect 2469 365 3445 367
rect 1477 316 1911 317
rect 1477 270 1836 316
rect 1882 270 1911 316
rect 1007 152 1053 215
rect 1477 153 1523 270
rect 2469 244 2515 365
rect 3496 312 3563 472
rect 2196 198 2209 244
rect 2255 198 2515 244
rect 2605 248 3563 312
rect 2605 192 2667 248
rect 1262 152 1523 153
rect 38 106 49 152
rect 95 106 106 152
rect 167 106 273 152
rect 319 106 330 152
rect 486 106 497 152
rect 543 106 554 152
rect 710 106 721 152
rect 767 106 1053 152
rect 1118 106 1129 152
rect 1175 106 1186 152
rect 1262 106 1273 152
rect 1319 106 1523 152
rect 1670 152 1738 155
rect 1670 106 1681 152
rect 1727 106 1738 152
rect 1912 106 1941 152
rect 1987 106 2477 152
rect 2523 106 2536 152
rect 2605 146 2621 192
rect 3053 192 3115 248
rect 2605 120 2667 146
rect 2845 152 2891 170
rect 3053 146 3069 192
rect 3501 191 3563 248
rect 3053 120 3115 146
rect 3293 155 3339 168
rect 38 60 106 106
rect 486 60 554 106
rect 1118 60 1186 106
rect 1670 60 1738 106
rect 2845 60 2891 106
rect 3501 145 3517 191
rect 3501 120 3563 145
rect 3293 60 3339 109
rect 0 -60 3696 60
<< labels >>
flabel metal1 s 1582 364 2120 423 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 3696 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2845 168 2891 170 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 3474 663 3563 665 0 FreeSans 400 0 0 0 Z
port 4 nsew default output
flabel metal1 s 376 253 872 307 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 173 491 420 542 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 173 445 775 491 1 A2
port 2 nsew default input
rlabel metal1 s 729 419 775 445 1 A2
port 2 nsew default input
rlabel metal1 s 173 419 221 445 1 A2
port 2 nsew default input
rlabel metal1 s 729 364 979 419 1 A2
port 2 nsew default input
rlabel metal1 s 173 364 221 419 1 A2
port 2 nsew default input
rlabel metal1 s 923 358 979 364 1 A2
port 2 nsew default input
rlabel metal1 s 173 358 221 364 1 A2
port 2 nsew default input
rlabel metal1 s 923 320 1072 358 1 A2
port 2 nsew default input
rlabel metal1 s 173 320 221 358 1 A2
port 2 nsew default input
rlabel metal1 s 923 312 1072 320 1 A2
port 2 nsew default input
rlabel metal1 s 3474 536 3563 663 1 Z
port 4 nsew default output
rlabel metal1 s 3053 536 3138 663 1 Z
port 4 nsew default output
rlabel metal1 s 2605 536 2701 663 1 Z
port 4 nsew default output
rlabel metal1 s 2605 472 3563 536 1 Z
port 4 nsew default output
rlabel metal1 s 3496 312 3563 472 1 Z
port 4 nsew default output
rlabel metal1 s 2605 248 3563 312 1 Z
port 4 nsew default output
rlabel metal1 s 3501 120 3563 248 1 Z
port 4 nsew default output
rlabel metal1 s 3053 120 3115 248 1 Z
port 4 nsew default output
rlabel metal1 s 2605 120 2667 248 1 Z
port 4 nsew default output
rlabel metal1 s 3283 657 3329 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2845 657 2891 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2446 657 2514 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1714 657 1782 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1273 657 1319 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 657 534 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3283 588 3329 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2845 588 2891 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1714 588 1782 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1273 588 1319 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 588 534 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1714 561 1782 588 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1273 561 1319 588 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 561 534 588 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1273 537 1319 561 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 537 534 561 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1273 497 1319 537 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3293 155 3339 168 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2845 155 2891 168 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3293 152 3339 155 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2845 152 2891 155 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1670 152 1738 155 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3293 60 3339 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2845 60 2891 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1670 60 1738 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1118 60 1186 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3696 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3696 784
string GDS_END 392658
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 384626
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
