magic
tech gf180mcuA
timestamp 1752776960
<< properties >>
string gencell npn_00p54x10p00_0
string library gf180mcu
string parameter m=1
<< end >>
