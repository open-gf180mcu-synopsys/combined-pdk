magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 565 390 635
rect 140 360 165 565
rect 225 390 250 530
rect 215 388 265 390
rect 215 362 227 388
rect 253 362 265 388
rect 215 360 265 362
rect 310 360 335 565
rect 105 258 155 260
rect 105 232 117 258
rect 143 232 155 258
rect 105 230 155 232
rect 140 70 165 190
rect 225 105 250 360
rect 310 70 335 190
rect 0 0 390 70
<< via1 >>
rect 227 362 253 388
rect 117 232 143 258
<< obsm1 >>
rect 55 335 80 530
rect 55 305 200 335
rect 55 105 80 305
<< metal2 >>
rect 215 388 265 395
rect 215 362 227 388
rect 253 362 265 388
rect 215 355 265 362
rect 110 260 150 265
rect 105 258 155 260
rect 105 232 117 258
rect 143 232 155 258
rect 105 230 155 232
rect 110 225 150 230
<< labels >>
rlabel metal1 s 140 360 165 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 310 360 335 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 565 390 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 140 0 165 190 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 310 0 335 190 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 0 390 70 6 VSS
port 4 nsew ground bidirectional abutment
rlabel via1 s 117 232 143 258 6 A
port 1 nsew signal input
rlabel metal2 s 110 225 150 265 6 A
port 1 nsew signal input
rlabel metal2 s 105 230 155 260 6 A
port 1 nsew signal input
rlabel metal1 s 105 230 155 260 6 A
port 1 nsew signal input
rlabel via1 s 227 362 253 388 6 Y
port 2 nsew signal output
rlabel metal2 s 215 355 265 395 6 Y
port 2 nsew signal output
rlabel metal1 s 225 105 250 530 6 Y
port 2 nsew signal output
rlabel metal1 s 215 360 265 390 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 390 635
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 104864
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 99840
<< end >>
