magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< isosubstrate >>
rect -83 -83 5981 8547
<< nwell >>
rect -83 6391 5981 8547
rect 454 3720 5444 5844
rect -83 2617 5981 3173
rect -83 473 473 2617
rect 5425 473 5981 2617
rect -83 -83 5981 473
<< psubdiff >>
rect 0 6305 5898 6327
rect 0 3259 22 6305
rect 368 5959 476 6305
rect 5422 5959 5530 6305
rect 368 5937 5530 5959
rect 368 3627 390 5937
rect 5508 3627 5530 5937
rect 368 3605 5530 3627
rect 368 3259 476 3605
rect 5422 3259 5530 3605
rect 5876 3259 5898 6305
rect 0 3237 5898 3259
rect 537 2502 5361 2524
rect 537 2456 576 2502
rect 5322 2456 5361 2502
rect 537 2348 5361 2456
rect 537 2320 858 2348
rect 537 770 559 2320
rect 605 1710 713 2320
rect 759 2302 858 2320
rect 5040 2320 5361 2348
rect 5040 2302 5139 2320
rect 759 2280 5139 2302
rect 759 1744 781 2280
rect 5117 1744 5139 2280
rect 759 1722 5139 1744
rect 759 1710 858 1722
rect 605 1676 858 1710
rect 5040 1710 5139 1722
rect 5185 1710 5293 2320
rect 5040 1676 5293 1710
rect 605 1568 5293 1676
rect 605 1522 717 1568
rect 5181 1522 5293 1568
rect 605 1414 5293 1522
rect 605 1386 858 1414
rect 605 776 713 1386
rect 759 1368 858 1386
rect 5040 1386 5293 1414
rect 5040 1368 5139 1386
rect 759 1346 5139 1368
rect 759 810 781 1346
rect 5117 810 5139 1346
rect 759 788 5139 810
rect 759 776 858 788
rect 605 770 858 776
rect 537 742 858 770
rect 5040 776 5139 788
rect 5185 776 5293 1386
rect 5040 770 5293 776
rect 5339 770 5361 2320
rect 5040 742 5361 770
rect 537 634 5361 742
rect 537 588 576 634
rect 5322 588 5361 634
rect 537 566 5361 588
<< nsubdiff >>
rect 0 8442 5898 8464
rect 0 6496 22 8442
rect 368 8096 476 8442
rect 5422 8096 5530 8442
rect 368 8074 5530 8096
rect 368 6864 390 8074
rect 5508 6864 5530 8074
rect 368 6842 5530 6864
rect 368 6496 476 6842
rect 5422 6496 5530 6842
rect 5876 6496 5898 8442
rect 0 6474 5898 6496
rect 537 5739 5361 5761
rect 537 5693 576 5739
rect 5322 5693 5361 5739
rect 537 5585 5361 5693
rect 537 5557 858 5585
rect 537 4007 559 5557
rect 605 4947 713 5557
rect 759 5539 858 5557
rect 5040 5557 5361 5585
rect 5040 5539 5139 5557
rect 759 5517 5139 5539
rect 759 4981 781 5517
rect 5117 4981 5139 5517
rect 759 4959 5139 4981
rect 759 4947 858 4959
rect 605 4913 858 4947
rect 5040 4947 5139 4959
rect 5185 4947 5293 5557
rect 5040 4913 5293 4947
rect 605 4805 5293 4913
rect 605 4759 717 4805
rect 5181 4759 5293 4805
rect 605 4651 5293 4759
rect 605 4623 858 4651
rect 605 4013 713 4623
rect 759 4605 858 4623
rect 5040 4623 5293 4651
rect 5040 4605 5139 4623
rect 759 4583 5139 4605
rect 759 4047 781 4583
rect 5117 4047 5139 4583
rect 759 4025 5139 4047
rect 759 4013 858 4025
rect 605 4007 858 4013
rect 537 3979 858 4007
rect 5040 4013 5139 4025
rect 5185 4013 5293 4623
rect 5040 4007 5293 4013
rect 5339 4007 5361 5557
rect 5040 3979 5361 4007
rect 537 3871 5361 3979
rect 537 3825 576 3871
rect 5322 3825 5361 3871
rect 537 3803 5361 3825
rect 0 3068 5898 3090
rect 0 22 22 3068
rect 368 2722 476 3068
rect 5422 2722 5530 3068
rect 368 2700 5530 2722
rect 368 390 390 2700
rect 5508 390 5530 2700
rect 368 368 5530 390
rect 368 22 476 368
rect 5422 22 5530 368
rect 5876 22 5898 3068
rect 0 0 5898 22
<< psubdiffcont >>
rect 22 3259 368 6305
rect 476 5959 5422 6305
rect 476 3259 5422 3605
rect 5530 3259 5876 6305
rect 576 2456 5322 2502
rect 559 770 605 2320
rect 713 1710 759 2320
rect 858 2302 5040 2348
rect 858 1676 5040 1722
rect 5139 1710 5185 2320
rect 717 1522 5181 1568
rect 713 776 759 1386
rect 858 1368 5040 1414
rect 858 742 5040 788
rect 5139 776 5185 1386
rect 5293 770 5339 2320
rect 576 588 5322 634
<< nsubdiffcont >>
rect 22 6496 368 8442
rect 476 8096 5422 8442
rect 476 6496 5422 6842
rect 5530 6496 5876 8442
rect 576 5693 5322 5739
rect 559 4007 605 5557
rect 713 4947 759 5557
rect 858 5539 5040 5585
rect 858 4913 5040 4959
rect 5139 4947 5185 5557
rect 717 4759 5181 4805
rect 713 4013 759 4623
rect 858 4605 5040 4651
rect 858 3979 5040 4025
rect 5139 4013 5185 4623
rect 5293 4007 5339 5557
rect 576 3825 5322 3871
rect 22 22 368 3068
rect 476 2722 5422 3068
rect 476 22 5422 368
rect 5530 22 5876 3068
<< polysilicon >>
rect 1769 7838 2269 7851
rect 1769 7792 1782 7838
rect 1828 7792 1889 7838
rect 1935 7792 1996 7838
rect 2042 7792 2103 7838
rect 2149 7792 2210 7838
rect 2256 7792 2269 7838
rect 1769 7749 2269 7792
rect 1769 7146 2269 7189
rect 1769 7100 1782 7146
rect 1828 7100 1889 7146
rect 1935 7100 1996 7146
rect 2042 7100 2103 7146
rect 2149 7100 2210 7146
rect 2256 7100 2269 7146
rect 1769 7087 2269 7100
rect 2389 7838 2889 7851
rect 2389 7792 2402 7838
rect 2448 7792 2509 7838
rect 2555 7792 2616 7838
rect 2662 7792 2723 7838
rect 2769 7792 2830 7838
rect 2876 7792 2889 7838
rect 2389 7749 2889 7792
rect 2389 7146 2889 7189
rect 2389 7100 2402 7146
rect 2448 7100 2509 7146
rect 2555 7100 2616 7146
rect 2662 7100 2723 7146
rect 2769 7100 2830 7146
rect 2876 7100 2889 7146
rect 2389 7087 2889 7100
rect 3009 7838 3509 7851
rect 3009 7792 3022 7838
rect 3068 7792 3129 7838
rect 3175 7792 3236 7838
rect 3282 7792 3343 7838
rect 3389 7792 3450 7838
rect 3496 7792 3509 7838
rect 3009 7749 3509 7792
rect 3009 7146 3509 7189
rect 3009 7100 3022 7146
rect 3068 7100 3129 7146
rect 3175 7100 3236 7146
rect 3282 7100 3343 7146
rect 3389 7100 3450 7146
rect 3496 7100 3509 7146
rect 3009 7087 3509 7100
rect 3629 7838 4129 7851
rect 3629 7792 3642 7838
rect 3688 7792 3749 7838
rect 3795 7792 3856 7838
rect 3902 7792 3963 7838
rect 4009 7792 4070 7838
rect 4116 7792 4129 7838
rect 3629 7749 4129 7792
rect 3629 7146 4129 7189
rect 3629 7100 3642 7146
rect 3688 7100 3749 7146
rect 3795 7100 3856 7146
rect 3902 7100 3963 7146
rect 4009 7100 4070 7146
rect 4116 7100 4129 7146
rect 3629 7087 4129 7100
<< polycontact >>
rect 1782 7792 1828 7838
rect 1889 7792 1935 7838
rect 1996 7792 2042 7838
rect 2103 7792 2149 7838
rect 2210 7792 2256 7838
rect 1782 7100 1828 7146
rect 1889 7100 1935 7146
rect 1996 7100 2042 7146
rect 2103 7100 2149 7146
rect 2210 7100 2256 7146
rect 2402 7792 2448 7838
rect 2509 7792 2555 7838
rect 2616 7792 2662 7838
rect 2723 7792 2769 7838
rect 2830 7792 2876 7838
rect 2402 7100 2448 7146
rect 2509 7100 2555 7146
rect 2616 7100 2662 7146
rect 2723 7100 2769 7146
rect 2830 7100 2876 7146
rect 3022 7792 3068 7838
rect 3129 7792 3175 7838
rect 3236 7792 3282 7838
rect 3343 7792 3389 7838
rect 3450 7792 3496 7838
rect 3022 7100 3068 7146
rect 3129 7100 3175 7146
rect 3236 7100 3282 7146
rect 3343 7100 3389 7146
rect 3450 7100 3496 7146
rect 3642 7792 3688 7838
rect 3749 7792 3795 7838
rect 3856 7792 3902 7838
rect 3963 7792 4009 7838
rect 4070 7792 4116 7838
rect 3642 7100 3688 7146
rect 3749 7100 3795 7146
rect 3856 7100 3902 7146
rect 3963 7100 4009 7146
rect 4070 7100 4116 7146
<< ppolyres >>
rect 1769 7189 2269 7749
rect 2389 7189 2889 7749
rect 3009 7189 3509 7749
rect 3629 7189 4129 7749
<< mvpdiode >>
rect 949 5336 4949 5349
rect 949 5290 962 5336
rect 4936 5290 4949 5336
rect 949 5208 4949 5290
rect 949 5162 962 5208
rect 4936 5162 4949 5208
rect 949 5149 4949 5162
rect 949 4402 4949 4415
rect 949 4356 962 4402
rect 4936 4356 4949 4402
rect 949 4274 4949 4356
rect 949 4228 962 4274
rect 4936 4228 4949 4274
rect 949 4215 4949 4228
<< mvndiode >>
rect 949 2099 4949 2112
rect 949 2053 962 2099
rect 4936 2053 4949 2099
rect 949 1971 4949 2053
rect 949 1925 962 1971
rect 4936 1925 4949 1971
rect 949 1912 4949 1925
rect 949 1165 4949 1178
rect 949 1119 962 1165
rect 4936 1119 4949 1165
rect 949 1037 4949 1119
rect 949 991 962 1037
rect 4936 991 4949 1037
rect 949 978 4949 991
<< mvpdiodec >>
rect 962 5290 4936 5336
rect 962 5162 4936 5208
rect 962 4356 4936 4402
rect 962 4228 4936 4274
<< mvndiodec >>
rect 962 2053 4936 2099
rect 962 1925 4936 1971
rect 962 1119 4936 1165
rect 962 991 4936 1037
<< metal1 >>
rect 11 8442 5887 8453
rect 11 6496 22 8442
rect 368 8403 476 8442
rect 5422 8403 5530 8442
rect 368 8351 466 8403
rect 5432 8351 5530 8403
rect 368 8295 476 8351
rect 5422 8295 5530 8351
rect 368 8243 466 8295
rect 5432 8243 5530 8295
rect 368 8187 476 8243
rect 5422 8187 5530 8243
rect 368 8135 466 8187
rect 5432 8135 5530 8187
rect 368 8096 476 8135
rect 5422 8096 5530 8135
rect 368 8085 5530 8096
rect 368 6853 379 8085
rect 1766 7949 4130 7961
rect 1766 7793 1778 7949
rect 4118 7793 4130 7949
rect 1766 7792 1782 7793
rect 1828 7792 1889 7793
rect 1935 7792 1996 7793
rect 2042 7792 2103 7793
rect 2149 7792 2210 7793
rect 2256 7792 2402 7793
rect 2448 7792 2509 7793
rect 2555 7792 2616 7793
rect 2662 7792 2723 7793
rect 2769 7792 2830 7793
rect 2876 7792 3022 7793
rect 3068 7792 3129 7793
rect 3175 7792 3236 7793
rect 3282 7792 3343 7793
rect 3389 7792 3450 7793
rect 3496 7792 3642 7793
rect 3688 7792 3749 7793
rect 3795 7792 3856 7793
rect 3902 7792 3963 7793
rect 4009 7792 4070 7793
rect 4116 7792 4130 7793
rect 1766 7781 4130 7792
rect 1766 7146 4130 7157
rect 1766 7145 1782 7146
rect 1828 7145 1889 7146
rect 1935 7145 1996 7146
rect 2042 7145 2103 7146
rect 2149 7145 2210 7146
rect 2256 7145 2402 7146
rect 2448 7145 2509 7146
rect 2555 7145 2616 7146
rect 2662 7145 2723 7146
rect 2769 7145 2830 7146
rect 2876 7145 3022 7146
rect 3068 7145 3129 7146
rect 3175 7145 3236 7146
rect 3282 7145 3343 7146
rect 3389 7145 3450 7146
rect 3496 7145 3642 7146
rect 3688 7145 3749 7146
rect 3795 7145 3856 7146
rect 3902 7145 3963 7146
rect 4009 7145 4070 7146
rect 4116 7145 4130 7146
rect 1766 6989 1778 7145
rect 4118 6989 4130 7145
rect 1766 6977 4130 6989
rect 5519 6853 5530 8085
rect 368 6842 5530 6853
rect 368 6496 476 6842
rect 5422 6496 5530 6842
rect 5876 6496 5887 8442
rect 11 6485 5887 6496
rect 11 6305 5887 6316
rect 11 3259 22 6305
rect 368 5959 476 6305
rect 5422 5959 5530 6305
rect 368 5948 5530 5959
rect 368 3616 379 5948
rect 548 5739 5350 5750
rect 548 5693 576 5739
rect 5322 5693 5350 5739
rect 548 5656 579 5693
rect 631 5656 687 5693
rect 739 5656 1496 5693
rect 548 5600 1496 5656
rect 548 5557 579 5600
rect 548 4007 559 5557
rect 631 5548 687 5600
rect 739 5585 1496 5600
rect 1860 5585 2508 5693
rect 2872 5585 3026 5693
rect 3390 5585 4038 5693
rect 4402 5656 5159 5693
rect 5211 5656 5267 5693
rect 5319 5656 5350 5693
rect 4402 5600 5350 5656
rect 4402 5585 5159 5600
rect 739 5557 858 5585
rect 605 5492 713 5548
rect 759 5539 858 5557
rect 5040 5557 5159 5585
rect 5040 5539 5139 5557
rect 5211 5548 5267 5600
rect 5319 5557 5350 5600
rect 759 5528 5139 5539
rect 631 5440 687 5492
rect 605 5384 713 5440
rect 631 5332 687 5384
rect 605 5276 713 5332
rect 631 5224 687 5276
rect 605 5168 713 5224
rect 631 5116 687 5168
rect 605 5060 713 5116
rect 631 5008 687 5060
rect 605 4952 713 5008
rect 759 4970 770 5528
rect 949 5336 4949 5349
rect 949 5290 962 5336
rect 4936 5290 4949 5336
rect 949 5208 990 5290
rect 1354 5208 2002 5290
rect 2366 5208 3532 5290
rect 3896 5208 4544 5290
rect 4908 5208 4949 5290
rect 949 5162 962 5208
rect 4936 5162 4949 5208
rect 949 5149 4949 5162
rect 5128 4970 5139 5528
rect 5185 5492 5293 5548
rect 5211 5440 5267 5492
rect 5185 5384 5293 5440
rect 5211 5332 5267 5384
rect 5185 5276 5293 5332
rect 5211 5224 5267 5276
rect 5185 5168 5293 5224
rect 5211 5116 5267 5168
rect 5185 5060 5293 5116
rect 5211 5008 5267 5060
rect 759 4959 5139 4970
rect 631 4900 687 4952
rect 759 4947 858 4959
rect 739 4913 858 4947
rect 5040 4947 5139 4959
rect 5185 4952 5293 5008
rect 5040 4913 5159 4947
rect 739 4912 5159 4913
rect 739 4900 1496 4912
rect 605 4805 1496 4900
rect 1860 4805 2508 4912
rect 2872 4805 3026 4912
rect 3390 4805 4038 4912
rect 4402 4900 5159 4912
rect 5211 4900 5267 4952
rect 4402 4805 5293 4900
rect 605 4759 717 4805
rect 5181 4759 5293 4805
rect 605 4652 1496 4759
rect 1860 4652 2508 4759
rect 2872 4652 3026 4759
rect 3390 4652 4038 4759
rect 4402 4652 5293 4759
rect 605 4651 5293 4652
rect 605 4623 858 4651
rect 605 4013 713 4623
rect 759 4605 858 4623
rect 5040 4623 5293 4651
rect 5040 4605 5139 4623
rect 759 4594 5139 4605
rect 759 4036 770 4594
rect 949 4402 4949 4415
rect 949 4356 962 4402
rect 4936 4356 4949 4402
rect 949 4274 990 4356
rect 1354 4274 2002 4356
rect 2366 4274 3532 4356
rect 3896 4274 4544 4356
rect 4908 4274 4949 4356
rect 949 4228 962 4274
rect 4936 4228 4949 4274
rect 949 4215 4949 4228
rect 5128 4036 5139 4594
rect 759 4025 5139 4036
rect 759 4013 858 4025
rect 605 4007 858 4013
rect 548 3979 858 4007
rect 5040 4013 5139 4025
rect 5185 4013 5293 4623
rect 5040 4007 5293 4013
rect 5339 4007 5350 5557
rect 5040 3979 5350 4007
rect 548 3871 1496 3979
rect 1860 3871 2508 3979
rect 2872 3871 3026 3979
rect 3390 3871 4038 3979
rect 4402 3871 5350 3979
rect 548 3825 576 3871
rect 5322 3825 5350 3871
rect 548 3814 5350 3825
rect 5519 3616 5530 5948
rect 368 3605 5530 3616
rect 368 3259 476 3605
rect 5422 3259 5530 3605
rect 5876 3259 5887 6305
rect 11 3248 5887 3259
rect 11 3068 5887 3079
rect 11 22 22 3068
rect 368 2722 476 3068
rect 5422 2722 5530 3068
rect 368 2711 5530 2722
rect 368 379 379 2711
rect 548 2502 5350 2513
rect 548 2456 576 2502
rect 5322 2456 5350 2502
rect 548 2348 1496 2456
rect 1860 2348 2556 2456
rect 2712 2348 3187 2456
rect 3343 2348 4038 2456
rect 4402 2348 5350 2456
rect 548 2320 858 2348
rect 548 770 559 2320
rect 605 1710 713 2320
rect 759 2302 858 2320
rect 5040 2320 5350 2348
rect 5040 2302 5139 2320
rect 759 2291 5139 2302
rect 759 1733 770 2291
rect 949 2099 4949 2112
rect 949 2053 962 2099
rect 4936 2053 4949 2099
rect 949 1971 990 2053
rect 1354 1971 2002 2053
rect 2366 1971 3532 2053
rect 3896 1971 4544 2053
rect 4908 1971 4949 2053
rect 949 1925 962 1971
rect 4936 1925 4949 1971
rect 949 1912 4949 1925
rect 5128 1733 5139 2291
rect 759 1722 5139 1733
rect 759 1710 858 1722
rect 605 1676 858 1710
rect 5040 1710 5139 1722
rect 5185 1710 5293 2320
rect 5040 1676 5293 1710
rect 605 1675 5293 1676
rect 605 1568 1496 1675
rect 1860 1568 2554 1675
rect 2710 1568 3185 1675
rect 3341 1568 4038 1675
rect 4402 1568 5293 1675
rect 605 1522 717 1568
rect 5181 1522 5293 1568
rect 605 1416 1496 1522
rect 631 1364 687 1416
rect 739 1415 1496 1416
rect 1860 1415 2554 1522
rect 2710 1415 3185 1522
rect 3341 1415 4038 1522
rect 4402 1416 5293 1522
rect 4402 1415 5159 1416
rect 739 1414 5159 1415
rect 739 1386 858 1414
rect 759 1368 858 1386
rect 5040 1386 5159 1414
rect 5040 1368 5139 1386
rect 605 1308 713 1364
rect 759 1357 5139 1368
rect 5211 1364 5267 1416
rect 631 1256 687 1308
rect 605 1200 713 1256
rect 631 1148 687 1200
rect 605 1092 713 1148
rect 631 1040 687 1092
rect 605 984 713 1040
rect 631 932 687 984
rect 605 876 713 932
rect 631 824 687 876
rect 605 776 713 824
rect 759 799 770 1357
rect 949 1165 4949 1178
rect 949 1119 962 1165
rect 4936 1119 4949 1165
rect 949 1037 990 1119
rect 1354 1037 2002 1119
rect 2366 1037 3532 1119
rect 3896 1037 4544 1119
rect 4908 1037 4949 1119
rect 949 991 962 1037
rect 4936 991 4949 1037
rect 949 978 4949 991
rect 5128 799 5139 1357
rect 5185 1308 5293 1364
rect 5211 1256 5267 1308
rect 5185 1200 5293 1256
rect 5211 1148 5267 1200
rect 5185 1092 5293 1148
rect 5211 1040 5267 1092
rect 5185 984 5293 1040
rect 5211 932 5267 984
rect 5185 876 5293 932
rect 5211 824 5267 876
rect 759 788 5139 799
rect 759 776 858 788
rect 605 770 858 776
rect 548 768 858 770
rect 5040 776 5139 788
rect 5185 776 5293 824
rect 5040 770 5293 776
rect 5339 770 5350 2320
rect 5040 768 5350 770
rect 548 716 579 768
rect 631 716 687 768
rect 739 716 817 768
rect 869 716 925 742
rect 977 716 1033 742
rect 1085 716 1141 742
rect 1193 716 1249 742
rect 1301 716 1357 742
rect 1409 716 1465 742
rect 1517 716 1573 742
rect 1625 716 1681 742
rect 1733 716 1789 742
rect 1841 716 1897 742
rect 1949 716 2005 742
rect 2057 716 2113 742
rect 2165 716 2221 742
rect 2273 716 2329 742
rect 2381 716 2437 742
rect 2489 716 2545 742
rect 2597 716 2653 742
rect 2705 716 3193 742
rect 3245 716 3301 742
rect 3353 716 3409 742
rect 3461 716 3517 742
rect 3569 716 3625 742
rect 3677 716 3733 742
rect 3785 716 3841 742
rect 3893 716 3949 742
rect 4001 716 4057 742
rect 4109 716 4165 742
rect 4217 716 4273 742
rect 4325 716 4381 742
rect 4433 716 4489 742
rect 4541 716 4597 742
rect 4649 716 4705 742
rect 4757 716 4813 742
rect 4865 716 4921 742
rect 4973 716 5029 742
rect 5081 716 5159 768
rect 5211 716 5267 768
rect 5319 716 5350 768
rect 548 660 5350 716
rect 548 634 579 660
rect 631 634 687 660
rect 739 634 817 660
rect 869 634 925 660
rect 977 634 1033 660
rect 1085 634 1141 660
rect 1193 634 1249 660
rect 1301 634 1357 660
rect 1409 634 1465 660
rect 1517 634 1573 660
rect 1625 634 1681 660
rect 1733 634 1789 660
rect 1841 634 1897 660
rect 1949 634 2005 660
rect 2057 634 2113 660
rect 2165 634 2221 660
rect 2273 634 2329 660
rect 2381 634 2437 660
rect 2489 634 2545 660
rect 2597 634 2653 660
rect 2705 634 3193 660
rect 3245 634 3301 660
rect 3353 634 3409 660
rect 3461 634 3517 660
rect 3569 634 3625 660
rect 3677 634 3733 660
rect 3785 634 3841 660
rect 3893 634 3949 660
rect 4001 634 4057 660
rect 4109 634 4165 660
rect 4217 634 4273 660
rect 4325 634 4381 660
rect 4433 634 4489 660
rect 4541 634 4597 660
rect 4649 634 4705 660
rect 4757 634 4813 660
rect 4865 634 4921 660
rect 4973 634 5029 660
rect 5081 634 5159 660
rect 5211 634 5267 660
rect 5319 634 5350 660
rect 548 588 576 634
rect 5322 588 5350 634
rect 548 577 5350 588
rect 5519 379 5530 2711
rect 368 368 5530 379
rect 368 22 476 368
rect 5422 22 5530 368
rect 5876 22 5887 3068
rect 11 11 5887 22
<< via1 >>
rect 61 8361 113 8413
rect 169 8361 221 8413
rect 277 8361 329 8413
rect 466 8351 476 8403
rect 476 8351 518 8403
rect 574 8351 626 8403
rect 682 8351 734 8403
rect 790 8351 842 8403
rect 898 8351 950 8403
rect 1006 8351 1058 8403
rect 1114 8351 1166 8403
rect 1222 8351 1274 8403
rect 1330 8351 1382 8403
rect 1438 8351 1490 8403
rect 1546 8351 1598 8403
rect 1654 8351 1706 8403
rect 1762 8351 1814 8403
rect 1870 8351 1922 8403
rect 1978 8351 2030 8403
rect 2086 8351 2138 8403
rect 2194 8351 2246 8403
rect 2302 8351 2354 8403
rect 2410 8351 2462 8403
rect 2518 8351 2570 8403
rect 3328 8351 3380 8403
rect 3436 8351 3488 8403
rect 3544 8351 3596 8403
rect 3652 8351 3704 8403
rect 3760 8351 3812 8403
rect 3868 8351 3920 8403
rect 3976 8351 4028 8403
rect 4084 8351 4136 8403
rect 4192 8351 4244 8403
rect 4300 8351 4352 8403
rect 4408 8351 4460 8403
rect 4516 8351 4568 8403
rect 4624 8351 4676 8403
rect 4732 8351 4784 8403
rect 4840 8351 4892 8403
rect 4948 8351 5000 8403
rect 5056 8351 5108 8403
rect 5164 8351 5216 8403
rect 5272 8351 5324 8403
rect 5380 8351 5422 8403
rect 5422 8351 5432 8403
rect 5569 8361 5621 8413
rect 5677 8361 5729 8413
rect 5785 8361 5837 8413
rect 61 8253 113 8305
rect 169 8253 221 8305
rect 277 8253 329 8305
rect 466 8243 476 8295
rect 476 8243 518 8295
rect 574 8243 626 8295
rect 682 8243 734 8295
rect 790 8243 842 8295
rect 898 8243 950 8295
rect 1006 8243 1058 8295
rect 1114 8243 1166 8295
rect 1222 8243 1274 8295
rect 1330 8243 1382 8295
rect 1438 8243 1490 8295
rect 1546 8243 1598 8295
rect 1654 8243 1706 8295
rect 1762 8243 1814 8295
rect 1870 8243 1922 8295
rect 1978 8243 2030 8295
rect 2086 8243 2138 8295
rect 2194 8243 2246 8295
rect 2302 8243 2354 8295
rect 2410 8243 2462 8295
rect 2518 8243 2570 8295
rect 3328 8243 3380 8295
rect 3436 8243 3488 8295
rect 3544 8243 3596 8295
rect 3652 8243 3704 8295
rect 3760 8243 3812 8295
rect 3868 8243 3920 8295
rect 3976 8243 4028 8295
rect 4084 8243 4136 8295
rect 4192 8243 4244 8295
rect 4300 8243 4352 8295
rect 4408 8243 4460 8295
rect 4516 8243 4568 8295
rect 4624 8243 4676 8295
rect 4732 8243 4784 8295
rect 4840 8243 4892 8295
rect 4948 8243 5000 8295
rect 5056 8243 5108 8295
rect 5164 8243 5216 8295
rect 5272 8243 5324 8295
rect 5380 8243 5422 8295
rect 5422 8243 5432 8295
rect 5569 8253 5621 8305
rect 5677 8253 5729 8305
rect 5785 8253 5837 8305
rect 61 8145 113 8197
rect 169 8145 221 8197
rect 277 8145 329 8197
rect 466 8135 476 8187
rect 476 8135 518 8187
rect 574 8135 626 8187
rect 682 8135 734 8187
rect 790 8135 842 8187
rect 898 8135 950 8187
rect 1006 8135 1058 8187
rect 1114 8135 1166 8187
rect 1222 8135 1274 8187
rect 1330 8135 1382 8187
rect 1438 8135 1490 8187
rect 1546 8135 1598 8187
rect 1654 8135 1706 8187
rect 1762 8135 1814 8187
rect 1870 8135 1922 8187
rect 1978 8135 2030 8187
rect 2086 8135 2138 8187
rect 2194 8135 2246 8187
rect 2302 8135 2354 8187
rect 2410 8135 2462 8187
rect 2518 8135 2570 8187
rect 3328 8135 3380 8187
rect 3436 8135 3488 8187
rect 3544 8135 3596 8187
rect 3652 8135 3704 8187
rect 3760 8135 3812 8187
rect 3868 8135 3920 8187
rect 3976 8135 4028 8187
rect 4084 8135 4136 8187
rect 4192 8135 4244 8187
rect 4300 8135 4352 8187
rect 4408 8135 4460 8187
rect 4516 8135 4568 8187
rect 4624 8135 4676 8187
rect 4732 8135 4784 8187
rect 4840 8135 4892 8187
rect 4948 8135 5000 8187
rect 5056 8135 5108 8187
rect 5164 8135 5216 8187
rect 5272 8135 5324 8187
rect 5380 8135 5422 8187
rect 5422 8135 5432 8187
rect 5569 8145 5621 8197
rect 5677 8145 5729 8197
rect 5785 8145 5837 8197
rect 61 8037 113 8089
rect 169 8037 221 8089
rect 277 8037 329 8089
rect 61 7929 113 7981
rect 169 7929 221 7981
rect 277 7929 329 7981
rect 61 7821 113 7873
rect 169 7821 221 7873
rect 277 7821 329 7873
rect 61 7713 113 7765
rect 169 7713 221 7765
rect 277 7713 329 7765
rect 61 7605 113 7657
rect 169 7605 221 7657
rect 277 7605 329 7657
rect 61 7497 113 7549
rect 169 7497 221 7549
rect 277 7497 329 7549
rect 61 7389 113 7441
rect 169 7389 221 7441
rect 277 7389 329 7441
rect 61 7281 113 7333
rect 169 7281 221 7333
rect 277 7281 329 7333
rect 61 7173 113 7225
rect 169 7173 221 7225
rect 277 7173 329 7225
rect 61 7065 113 7117
rect 169 7065 221 7117
rect 277 7065 329 7117
rect 61 6957 113 7009
rect 169 6957 221 7009
rect 277 6957 329 7009
rect 61 6849 113 6901
rect 169 6849 221 6901
rect 277 6849 329 6901
rect 1778 7838 4118 7949
rect 1778 7793 1782 7838
rect 1782 7793 1828 7838
rect 1828 7793 1889 7838
rect 1889 7793 1935 7838
rect 1935 7793 1996 7838
rect 1996 7793 2042 7838
rect 2042 7793 2103 7838
rect 2103 7793 2149 7838
rect 2149 7793 2210 7838
rect 2210 7793 2256 7838
rect 2256 7793 2402 7838
rect 2402 7793 2448 7838
rect 2448 7793 2509 7838
rect 2509 7793 2555 7838
rect 2555 7793 2616 7838
rect 2616 7793 2662 7838
rect 2662 7793 2723 7838
rect 2723 7793 2769 7838
rect 2769 7793 2830 7838
rect 2830 7793 2876 7838
rect 2876 7793 3022 7838
rect 3022 7793 3068 7838
rect 3068 7793 3129 7838
rect 3129 7793 3175 7838
rect 3175 7793 3236 7838
rect 3236 7793 3282 7838
rect 3282 7793 3343 7838
rect 3343 7793 3389 7838
rect 3389 7793 3450 7838
rect 3450 7793 3496 7838
rect 3496 7793 3642 7838
rect 3642 7793 3688 7838
rect 3688 7793 3749 7838
rect 3749 7793 3795 7838
rect 3795 7793 3856 7838
rect 3856 7793 3902 7838
rect 3902 7793 3963 7838
rect 3963 7793 4009 7838
rect 4009 7793 4070 7838
rect 4070 7793 4116 7838
rect 4116 7793 4118 7838
rect 1778 7100 1782 7145
rect 1782 7100 1828 7145
rect 1828 7100 1889 7145
rect 1889 7100 1935 7145
rect 1935 7100 1996 7145
rect 1996 7100 2042 7145
rect 2042 7100 2103 7145
rect 2103 7100 2149 7145
rect 2149 7100 2210 7145
rect 2210 7100 2256 7145
rect 2256 7100 2402 7145
rect 2402 7100 2448 7145
rect 2448 7100 2509 7145
rect 2509 7100 2555 7145
rect 2555 7100 2616 7145
rect 2616 7100 2662 7145
rect 2662 7100 2723 7145
rect 2723 7100 2769 7145
rect 2769 7100 2830 7145
rect 2830 7100 2876 7145
rect 2876 7100 3022 7145
rect 3022 7100 3068 7145
rect 3068 7100 3129 7145
rect 3129 7100 3175 7145
rect 3175 7100 3236 7145
rect 3236 7100 3282 7145
rect 3282 7100 3343 7145
rect 3343 7100 3389 7145
rect 3389 7100 3450 7145
rect 3450 7100 3496 7145
rect 3496 7100 3642 7145
rect 3642 7100 3688 7145
rect 3688 7100 3749 7145
rect 3749 7100 3795 7145
rect 3795 7100 3856 7145
rect 3856 7100 3902 7145
rect 3902 7100 3963 7145
rect 3963 7100 4009 7145
rect 4009 7100 4070 7145
rect 4070 7100 4116 7145
rect 4116 7100 4118 7145
rect 1778 6989 4118 7100
rect 5569 8037 5621 8089
rect 5677 8037 5729 8089
rect 5785 8037 5837 8089
rect 5569 7929 5621 7981
rect 5677 7929 5729 7981
rect 5785 7929 5837 7981
rect 5569 7821 5621 7873
rect 5677 7821 5729 7873
rect 5785 7821 5837 7873
rect 5569 7713 5621 7765
rect 5677 7713 5729 7765
rect 5785 7713 5837 7765
rect 5569 7605 5621 7657
rect 5677 7605 5729 7657
rect 5785 7605 5837 7657
rect 5569 7497 5621 7549
rect 5677 7497 5729 7549
rect 5785 7497 5837 7549
rect 5569 7389 5621 7441
rect 5677 7389 5729 7441
rect 5785 7389 5837 7441
rect 5569 7281 5621 7333
rect 5677 7281 5729 7333
rect 5785 7281 5837 7333
rect 5569 7173 5621 7225
rect 5677 7173 5729 7225
rect 5785 7173 5837 7225
rect 5569 7065 5621 7117
rect 5677 7065 5729 7117
rect 5785 7065 5837 7117
rect 5569 6957 5621 7009
rect 5677 6957 5729 7009
rect 5785 6957 5837 7009
rect 5569 6849 5621 6901
rect 5677 6849 5729 6901
rect 5785 6849 5837 6901
rect 61 6741 113 6793
rect 169 6741 221 6793
rect 277 6741 329 6793
rect 61 6633 113 6685
rect 169 6633 221 6685
rect 277 6633 329 6685
rect 61 6525 113 6577
rect 169 6525 221 6577
rect 277 6525 329 6577
rect 5569 6741 5621 6793
rect 5677 6741 5729 6793
rect 5785 6741 5837 6793
rect 5569 6633 5621 6685
rect 5677 6633 5729 6685
rect 5785 6633 5837 6685
rect 5569 6525 5621 6577
rect 5677 6525 5729 6577
rect 5785 6525 5837 6577
rect 61 4559 113 4611
rect 169 4559 221 4611
rect 277 4559 329 4611
rect 61 4451 113 4503
rect 169 4451 221 4503
rect 277 4451 329 4503
rect 61 4343 113 4395
rect 169 4343 221 4395
rect 277 4343 329 4395
rect 61 4235 113 4287
rect 169 4235 221 4287
rect 277 4235 329 4287
rect 61 4127 113 4179
rect 169 4127 221 4179
rect 277 4127 329 4179
rect 61 4019 113 4071
rect 169 4019 221 4071
rect 277 4019 329 4071
rect 61 3911 113 3963
rect 169 3911 221 3963
rect 277 3911 329 3963
rect 61 3803 113 3855
rect 169 3803 221 3855
rect 277 3803 329 3855
rect 61 3695 113 3747
rect 169 3695 221 3747
rect 277 3695 329 3747
rect 61 3587 113 3639
rect 169 3587 221 3639
rect 277 3587 329 3639
rect 579 5693 631 5708
rect 687 5693 739 5708
rect 1496 5693 1860 5717
rect 2508 5693 2872 5717
rect 3026 5693 3390 5717
rect 4038 5693 4402 5717
rect 5159 5693 5211 5708
rect 5267 5693 5319 5708
rect 579 5656 631 5693
rect 687 5656 739 5693
rect 579 5557 631 5600
rect 579 5548 605 5557
rect 605 5548 631 5557
rect 687 5557 739 5600
rect 1496 5585 1860 5693
rect 2508 5585 2872 5693
rect 3026 5585 3390 5693
rect 4038 5585 4402 5693
rect 5159 5656 5211 5693
rect 5267 5656 5319 5693
rect 1496 5561 1860 5585
rect 2508 5561 2872 5585
rect 3026 5561 3390 5585
rect 4038 5561 4402 5585
rect 687 5548 713 5557
rect 713 5548 739 5557
rect 5159 5557 5211 5600
rect 5159 5548 5185 5557
rect 5185 5548 5211 5557
rect 5267 5557 5319 5600
rect 5267 5548 5293 5557
rect 5293 5548 5319 5557
rect 579 5440 605 5492
rect 605 5440 631 5492
rect 687 5440 713 5492
rect 713 5440 739 5492
rect 579 5332 605 5384
rect 605 5332 631 5384
rect 687 5332 713 5384
rect 713 5332 739 5384
rect 579 5224 605 5276
rect 605 5224 631 5276
rect 687 5224 713 5276
rect 713 5224 739 5276
rect 579 5116 605 5168
rect 605 5116 631 5168
rect 687 5116 713 5168
rect 713 5116 739 5168
rect 579 5008 605 5060
rect 605 5008 631 5060
rect 687 5008 713 5060
rect 713 5008 739 5060
rect 990 5290 1354 5327
rect 2002 5290 2366 5327
rect 3532 5290 3896 5327
rect 4544 5290 4908 5327
rect 990 5208 1354 5290
rect 2002 5208 2366 5290
rect 3532 5208 3896 5290
rect 4544 5208 4908 5290
rect 990 5171 1354 5208
rect 2002 5171 2366 5208
rect 3532 5171 3896 5208
rect 4544 5171 4908 5208
rect 5159 5440 5185 5492
rect 5185 5440 5211 5492
rect 5267 5440 5293 5492
rect 5293 5440 5319 5492
rect 5159 5332 5185 5384
rect 5185 5332 5211 5384
rect 5267 5332 5293 5384
rect 5293 5332 5319 5384
rect 5159 5224 5185 5276
rect 5185 5224 5211 5276
rect 5267 5224 5293 5276
rect 5293 5224 5319 5276
rect 5159 5116 5185 5168
rect 5185 5116 5211 5168
rect 5267 5116 5293 5168
rect 5293 5116 5319 5168
rect 5159 5008 5185 5060
rect 5185 5008 5211 5060
rect 5267 5008 5293 5060
rect 5293 5008 5319 5060
rect 579 4900 605 4952
rect 605 4900 631 4952
rect 687 4947 713 4952
rect 713 4947 739 4952
rect 687 4900 739 4947
rect 5159 4947 5185 4952
rect 5185 4947 5211 4952
rect 1496 4805 1860 4912
rect 2508 4805 2872 4912
rect 3026 4805 3390 4912
rect 4038 4805 4402 4912
rect 5159 4900 5211 4947
rect 5267 4900 5293 4952
rect 5293 4900 5319 4952
rect 1496 4759 1860 4805
rect 2508 4759 2872 4805
rect 3026 4759 3390 4805
rect 4038 4759 4402 4805
rect 1496 4652 1860 4759
rect 2508 4652 2872 4759
rect 3026 4652 3390 4759
rect 4038 4652 4402 4759
rect 990 4356 1354 4393
rect 2002 4356 2366 4393
rect 3532 4356 3896 4393
rect 4544 4356 4908 4393
rect 990 4274 1354 4356
rect 2002 4274 2366 4356
rect 3532 4274 3896 4356
rect 4544 4274 4908 4356
rect 990 4237 1354 4274
rect 2002 4237 2366 4274
rect 3532 4237 3896 4274
rect 4544 4237 4908 4274
rect 1496 3979 1860 4003
rect 2508 3979 2872 4003
rect 3026 3979 3390 4003
rect 4038 3979 4402 4003
rect 1496 3871 1860 3979
rect 2508 3871 2872 3979
rect 3026 3871 3390 3979
rect 4038 3871 4402 3979
rect 1496 3847 1860 3871
rect 2508 3847 2872 3871
rect 3026 3847 3390 3871
rect 4038 3847 4402 3871
rect 5569 4581 5621 4633
rect 5677 4581 5729 4633
rect 5785 4581 5837 4633
rect 5569 4473 5621 4525
rect 5677 4473 5729 4525
rect 5785 4473 5837 4525
rect 5569 4365 5621 4417
rect 5677 4365 5729 4417
rect 5785 4365 5837 4417
rect 5569 4257 5621 4309
rect 5677 4257 5729 4309
rect 5785 4257 5837 4309
rect 5569 4149 5621 4201
rect 5677 4149 5729 4201
rect 5785 4149 5837 4201
rect 5569 4041 5621 4093
rect 5677 4041 5729 4093
rect 5785 4041 5837 4093
rect 5569 3933 5621 3985
rect 5677 3933 5729 3985
rect 5785 3933 5837 3985
rect 5569 3825 5621 3877
rect 5677 3825 5729 3877
rect 5785 3825 5837 3877
rect 5569 3717 5621 3769
rect 5677 3717 5729 3769
rect 5785 3717 5837 3769
rect 5569 3609 5621 3661
rect 5677 3609 5729 3661
rect 5785 3609 5837 3661
rect 5569 3501 5621 3553
rect 5677 3501 5729 3553
rect 5785 3501 5837 3553
rect 5569 3393 5621 3445
rect 5677 3393 5729 3445
rect 5785 3393 5837 3445
rect 5569 3285 5621 3337
rect 5677 3285 5729 3337
rect 5785 3285 5837 3337
rect 61 2769 113 2821
rect 169 2769 221 2821
rect 277 2769 329 2821
rect 5569 2981 5621 3033
rect 5677 2981 5729 3033
rect 5785 2981 5837 3033
rect 5569 2873 5621 2925
rect 5677 2873 5729 2925
rect 5785 2873 5837 2925
rect 5569 2765 5621 2817
rect 5677 2765 5729 2817
rect 5785 2765 5837 2817
rect 61 2661 113 2713
rect 169 2661 221 2713
rect 277 2661 329 2713
rect 61 2553 113 2605
rect 169 2553 221 2605
rect 277 2553 329 2605
rect 61 2445 113 2497
rect 169 2445 221 2497
rect 277 2445 329 2497
rect 61 2337 113 2389
rect 169 2337 221 2389
rect 277 2337 329 2389
rect 61 2229 113 2281
rect 169 2229 221 2281
rect 277 2229 329 2281
rect 61 2121 113 2173
rect 169 2121 221 2173
rect 277 2121 329 2173
rect 61 2013 113 2065
rect 169 2013 221 2065
rect 277 2013 329 2065
rect 61 1905 113 1957
rect 169 1905 221 1957
rect 277 1905 329 1957
rect 61 1797 113 1849
rect 169 1797 221 1849
rect 277 1797 329 1849
rect 61 1689 113 1741
rect 169 1689 221 1741
rect 277 1689 329 1741
rect 1496 2456 1860 2480
rect 2556 2456 2712 2480
rect 3187 2456 3343 2480
rect 4038 2456 4402 2480
rect 1496 2348 1860 2456
rect 2556 2348 2712 2456
rect 3187 2348 3343 2456
rect 4038 2348 4402 2456
rect 1496 2324 1860 2348
rect 2556 2324 2712 2348
rect 3187 2324 3343 2348
rect 4038 2324 4402 2348
rect 990 2053 1354 2090
rect 2002 2053 2366 2090
rect 3532 2053 3896 2090
rect 4544 2053 4908 2090
rect 990 1971 1354 2053
rect 2002 1971 2366 2053
rect 3532 1971 3896 2053
rect 4544 1971 4908 2053
rect 990 1934 1354 1971
rect 2002 1934 2366 1971
rect 3532 1934 3896 1971
rect 4544 1934 4908 1971
rect 1496 1568 1860 1675
rect 2554 1568 2710 1675
rect 3185 1568 3341 1675
rect 4038 1568 4402 1675
rect 1496 1522 1860 1568
rect 2554 1522 2710 1568
rect 3185 1522 3341 1568
rect 4038 1522 4402 1568
rect 579 1364 605 1416
rect 605 1364 631 1416
rect 687 1386 739 1416
rect 1496 1415 1860 1522
rect 2554 1415 2710 1522
rect 3185 1415 3341 1522
rect 4038 1415 4402 1522
rect 687 1364 713 1386
rect 713 1364 739 1386
rect 5159 1386 5211 1416
rect 5159 1364 5185 1386
rect 5185 1364 5211 1386
rect 5267 1364 5293 1416
rect 5293 1364 5319 1416
rect 579 1256 605 1308
rect 605 1256 631 1308
rect 687 1256 713 1308
rect 713 1256 739 1308
rect 579 1148 605 1200
rect 605 1148 631 1200
rect 687 1148 713 1200
rect 713 1148 739 1200
rect 579 1040 605 1092
rect 605 1040 631 1092
rect 687 1040 713 1092
rect 713 1040 739 1092
rect 579 932 605 984
rect 605 932 631 984
rect 687 932 713 984
rect 713 932 739 984
rect 579 824 605 876
rect 605 824 631 876
rect 687 824 713 876
rect 713 824 739 876
rect 990 1119 1354 1156
rect 2002 1119 2366 1156
rect 3532 1119 3896 1156
rect 4544 1119 4908 1156
rect 990 1037 1354 1119
rect 2002 1037 2366 1119
rect 3532 1037 3896 1119
rect 4544 1037 4908 1119
rect 990 1000 1354 1037
rect 2002 1000 2366 1037
rect 3532 1000 3896 1037
rect 4544 1000 4908 1037
rect 5159 1256 5185 1308
rect 5185 1256 5211 1308
rect 5267 1256 5293 1308
rect 5293 1256 5319 1308
rect 5159 1148 5185 1200
rect 5185 1148 5211 1200
rect 5267 1148 5293 1200
rect 5293 1148 5319 1200
rect 5159 1040 5185 1092
rect 5185 1040 5211 1092
rect 5267 1040 5293 1092
rect 5293 1040 5319 1092
rect 5159 932 5185 984
rect 5185 932 5211 984
rect 5267 932 5293 984
rect 5293 932 5319 984
rect 5159 824 5185 876
rect 5185 824 5211 876
rect 5267 824 5293 876
rect 5293 824 5319 876
rect 579 716 631 768
rect 687 716 739 768
rect 817 742 858 768
rect 858 742 869 768
rect 925 742 977 768
rect 1033 742 1085 768
rect 1141 742 1193 768
rect 1249 742 1301 768
rect 1357 742 1409 768
rect 1465 742 1517 768
rect 1573 742 1625 768
rect 1681 742 1733 768
rect 1789 742 1841 768
rect 1897 742 1949 768
rect 2005 742 2057 768
rect 2113 742 2165 768
rect 2221 742 2273 768
rect 2329 742 2381 768
rect 2437 742 2489 768
rect 2545 742 2597 768
rect 2653 742 2705 768
rect 3193 742 3245 768
rect 3301 742 3353 768
rect 3409 742 3461 768
rect 3517 742 3569 768
rect 3625 742 3677 768
rect 3733 742 3785 768
rect 3841 742 3893 768
rect 3949 742 4001 768
rect 4057 742 4109 768
rect 4165 742 4217 768
rect 4273 742 4325 768
rect 4381 742 4433 768
rect 4489 742 4541 768
rect 4597 742 4649 768
rect 4705 742 4757 768
rect 4813 742 4865 768
rect 4921 742 4973 768
rect 5029 742 5040 768
rect 5040 742 5081 768
rect 817 716 869 742
rect 925 716 977 742
rect 1033 716 1085 742
rect 1141 716 1193 742
rect 1249 716 1301 742
rect 1357 716 1409 742
rect 1465 716 1517 742
rect 1573 716 1625 742
rect 1681 716 1733 742
rect 1789 716 1841 742
rect 1897 716 1949 742
rect 2005 716 2057 742
rect 2113 716 2165 742
rect 2221 716 2273 742
rect 2329 716 2381 742
rect 2437 716 2489 742
rect 2545 716 2597 742
rect 2653 716 2705 742
rect 3193 716 3245 742
rect 3301 716 3353 742
rect 3409 716 3461 742
rect 3517 716 3569 742
rect 3625 716 3677 742
rect 3733 716 3785 742
rect 3841 716 3893 742
rect 3949 716 4001 742
rect 4057 716 4109 742
rect 4165 716 4217 742
rect 4273 716 4325 742
rect 4381 716 4433 742
rect 4489 716 4541 742
rect 4597 716 4649 742
rect 4705 716 4757 742
rect 4813 716 4865 742
rect 4921 716 4973 742
rect 5029 716 5081 742
rect 5159 716 5211 768
rect 5267 716 5319 768
rect 579 634 631 660
rect 687 634 739 660
rect 817 634 869 660
rect 925 634 977 660
rect 1033 634 1085 660
rect 1141 634 1193 660
rect 1249 634 1301 660
rect 1357 634 1409 660
rect 1465 634 1517 660
rect 1573 634 1625 660
rect 1681 634 1733 660
rect 1789 634 1841 660
rect 1897 634 1949 660
rect 2005 634 2057 660
rect 2113 634 2165 660
rect 2221 634 2273 660
rect 2329 634 2381 660
rect 2437 634 2489 660
rect 2545 634 2597 660
rect 2653 634 2705 660
rect 3193 634 3245 660
rect 3301 634 3353 660
rect 3409 634 3461 660
rect 3517 634 3569 660
rect 3625 634 3677 660
rect 3733 634 3785 660
rect 3841 634 3893 660
rect 3949 634 4001 660
rect 4057 634 4109 660
rect 4165 634 4217 660
rect 4273 634 4325 660
rect 4381 634 4433 660
rect 4489 634 4541 660
rect 4597 634 4649 660
rect 4705 634 4757 660
rect 4813 634 4865 660
rect 4921 634 4973 660
rect 5029 634 5081 660
rect 5159 634 5211 660
rect 5267 634 5319 660
rect 579 608 631 634
rect 687 608 739 634
rect 817 608 869 634
rect 925 608 977 634
rect 1033 608 1085 634
rect 1141 608 1193 634
rect 1249 608 1301 634
rect 1357 608 1409 634
rect 1465 608 1517 634
rect 1573 608 1625 634
rect 1681 608 1733 634
rect 1789 608 1841 634
rect 1897 608 1949 634
rect 2005 608 2057 634
rect 2113 608 2165 634
rect 2221 608 2273 634
rect 2329 608 2381 634
rect 2437 608 2489 634
rect 2545 608 2597 634
rect 2653 608 2705 634
rect 3193 608 3245 634
rect 3301 608 3353 634
rect 3409 608 3461 634
rect 3517 608 3569 634
rect 3625 608 3677 634
rect 3733 608 3785 634
rect 3841 608 3893 634
rect 3949 608 4001 634
rect 4057 608 4109 634
rect 4165 608 4217 634
rect 4273 608 4325 634
rect 4381 608 4433 634
rect 4489 608 4541 634
rect 4597 608 4649 634
rect 4705 608 4757 634
rect 4813 608 4865 634
rect 4921 608 4973 634
rect 5029 608 5081 634
rect 5159 608 5211 634
rect 5267 608 5319 634
rect 5569 2657 5621 2709
rect 5677 2657 5729 2709
rect 5785 2657 5837 2709
rect 5569 2549 5621 2601
rect 5677 2549 5729 2601
rect 5785 2549 5837 2601
rect 5569 2441 5621 2493
rect 5677 2441 5729 2493
rect 5785 2441 5837 2493
rect 5569 2333 5621 2385
rect 5677 2333 5729 2385
rect 5785 2333 5837 2385
rect 5569 2225 5621 2277
rect 5677 2225 5729 2277
rect 5785 2225 5837 2277
rect 5569 2117 5621 2169
rect 5677 2117 5729 2169
rect 5785 2117 5837 2169
rect 5569 2009 5621 2061
rect 5677 2009 5729 2061
rect 5785 2009 5837 2061
rect 5569 1901 5621 1953
rect 5677 1901 5729 1953
rect 5785 1901 5837 1953
rect 5569 1793 5621 1845
rect 5677 1793 5729 1845
rect 5785 1793 5837 1845
rect 5569 1685 5621 1737
rect 5677 1685 5729 1737
rect 5785 1685 5837 1737
<< metal2 >>
rect 11 8439 2582 8453
rect 11 8383 25 8439
rect 81 8413 167 8439
rect 223 8413 309 8439
rect 113 8383 167 8413
rect 223 8383 277 8413
rect 365 8383 451 8439
rect 507 8403 593 8439
rect 649 8403 735 8439
rect 791 8403 877 8439
rect 933 8403 1019 8439
rect 1075 8403 1161 8439
rect 1217 8403 1303 8439
rect 1359 8403 1445 8439
rect 1501 8403 1587 8439
rect 1643 8403 1729 8439
rect 1785 8403 1871 8439
rect 1927 8403 2013 8439
rect 2069 8403 2155 8439
rect 2211 8403 2297 8439
rect 2353 8403 2439 8439
rect 2495 8403 2582 8439
rect 11 8361 61 8383
rect 113 8361 169 8383
rect 221 8361 277 8383
rect 329 8361 466 8383
rect 11 8351 466 8361
rect 518 8351 574 8403
rect 649 8383 682 8403
rect 626 8351 682 8383
rect 734 8383 735 8403
rect 842 8383 877 8403
rect 734 8351 790 8383
rect 842 8351 898 8383
rect 950 8351 1006 8403
rect 1075 8383 1114 8403
rect 1217 8383 1222 8403
rect 1058 8351 1114 8383
rect 1166 8351 1222 8383
rect 1274 8383 1303 8403
rect 1274 8351 1330 8383
rect 1382 8351 1438 8403
rect 1501 8383 1546 8403
rect 1643 8383 1654 8403
rect 1490 8351 1546 8383
rect 1598 8351 1654 8383
rect 1706 8383 1729 8403
rect 1706 8351 1762 8383
rect 1814 8351 1870 8403
rect 1927 8383 1978 8403
rect 2069 8383 2086 8403
rect 1922 8351 1978 8383
rect 2030 8351 2086 8383
rect 2138 8383 2155 8403
rect 2246 8383 2297 8403
rect 2138 8351 2194 8383
rect 2246 8351 2302 8383
rect 2354 8351 2410 8403
rect 2495 8383 2518 8403
rect 2462 8351 2518 8383
rect 2570 8351 2582 8403
rect 11 8305 2582 8351
rect 11 8297 61 8305
rect 113 8297 169 8305
rect 221 8297 277 8305
rect 329 8297 2582 8305
rect 11 8241 25 8297
rect 113 8253 167 8297
rect 223 8253 277 8297
rect 81 8241 167 8253
rect 223 8241 309 8253
rect 365 8241 451 8297
rect 507 8295 593 8297
rect 649 8295 735 8297
rect 791 8295 877 8297
rect 933 8295 1019 8297
rect 1075 8295 1161 8297
rect 1217 8295 1303 8297
rect 1359 8295 1445 8297
rect 1501 8295 1587 8297
rect 1643 8295 1729 8297
rect 1785 8295 1871 8297
rect 1927 8295 2013 8297
rect 2069 8295 2155 8297
rect 2211 8295 2297 8297
rect 2353 8295 2439 8297
rect 2495 8295 2582 8297
rect 518 8243 574 8295
rect 649 8243 682 8295
rect 734 8243 735 8295
rect 842 8243 877 8295
rect 950 8243 1006 8295
rect 1075 8243 1114 8295
rect 1217 8243 1222 8295
rect 1274 8243 1303 8295
rect 1382 8243 1438 8295
rect 1501 8243 1546 8295
rect 1643 8243 1654 8295
rect 1706 8243 1729 8295
rect 1814 8243 1870 8295
rect 1927 8243 1978 8295
rect 2069 8243 2086 8295
rect 2138 8243 2155 8295
rect 2246 8243 2297 8295
rect 2354 8243 2410 8295
rect 2495 8243 2518 8295
rect 2570 8243 2582 8295
rect 507 8241 593 8243
rect 649 8241 735 8243
rect 791 8241 877 8243
rect 933 8241 1019 8243
rect 1075 8241 1161 8243
rect 1217 8241 1303 8243
rect 1359 8241 1445 8243
rect 1501 8241 1587 8243
rect 1643 8241 1729 8243
rect 1785 8241 1871 8243
rect 1927 8241 2013 8243
rect 2069 8241 2155 8243
rect 2211 8241 2297 8243
rect 2353 8241 2439 8243
rect 2495 8241 2582 8243
rect 11 8197 2582 8241
rect 11 8155 61 8197
rect 113 8155 169 8197
rect 221 8155 277 8197
rect 329 8187 2582 8197
rect 329 8155 466 8187
rect 11 8099 25 8155
rect 113 8145 167 8155
rect 223 8145 277 8155
rect 81 8099 167 8145
rect 223 8099 309 8145
rect 365 8099 451 8155
rect 518 8135 574 8187
rect 626 8155 682 8187
rect 649 8135 682 8155
rect 734 8155 790 8187
rect 842 8155 898 8187
rect 734 8135 735 8155
rect 842 8135 877 8155
rect 950 8135 1006 8187
rect 1058 8155 1114 8187
rect 1166 8155 1222 8187
rect 1075 8135 1114 8155
rect 1217 8135 1222 8155
rect 1274 8155 1330 8187
rect 1274 8135 1303 8155
rect 1382 8135 1438 8187
rect 1490 8155 1546 8187
rect 1598 8155 1654 8187
rect 1501 8135 1546 8155
rect 1643 8135 1654 8155
rect 1706 8155 1762 8187
rect 1706 8135 1729 8155
rect 1814 8135 1870 8187
rect 1922 8155 1978 8187
rect 2030 8155 2086 8187
rect 1927 8135 1978 8155
rect 2069 8135 2086 8155
rect 2138 8155 2194 8187
rect 2246 8155 2302 8187
rect 2138 8135 2155 8155
rect 2246 8135 2297 8155
rect 2354 8135 2410 8187
rect 2462 8155 2518 8187
rect 2495 8135 2518 8155
rect 2570 8135 2582 8187
rect 507 8099 593 8135
rect 649 8099 735 8135
rect 791 8099 877 8135
rect 933 8099 1019 8135
rect 1075 8099 1161 8135
rect 1217 8099 1303 8135
rect 1359 8099 1445 8135
rect 1501 8099 1587 8135
rect 1643 8099 1729 8135
rect 1785 8099 1871 8135
rect 1927 8099 2013 8135
rect 2069 8099 2155 8135
rect 2211 8099 2297 8135
rect 2353 8099 2439 8135
rect 2495 8099 2582 8135
rect 11 8089 2582 8099
rect 11 8037 61 8089
rect 113 8037 169 8089
rect 221 8037 277 8089
rect 329 8085 2582 8089
rect 3316 8439 5887 8453
rect 3316 8403 3403 8439
rect 3459 8403 3545 8439
rect 3601 8403 3687 8439
rect 3743 8403 3829 8439
rect 3885 8403 3971 8439
rect 4027 8403 4113 8439
rect 4169 8403 4255 8439
rect 4311 8403 4397 8439
rect 4453 8403 4539 8439
rect 4595 8403 4681 8439
rect 4737 8403 4823 8439
rect 4879 8403 4965 8439
rect 5021 8403 5107 8439
rect 5163 8403 5249 8439
rect 5305 8403 5391 8439
rect 3316 8351 3328 8403
rect 3380 8383 3403 8403
rect 3380 8351 3436 8383
rect 3488 8351 3544 8403
rect 3601 8383 3652 8403
rect 3743 8383 3760 8403
rect 3596 8351 3652 8383
rect 3704 8351 3760 8383
rect 3812 8383 3829 8403
rect 3920 8383 3971 8403
rect 3812 8351 3868 8383
rect 3920 8351 3976 8383
rect 4028 8351 4084 8403
rect 4169 8383 4192 8403
rect 4136 8351 4192 8383
rect 4244 8383 4255 8403
rect 4352 8383 4397 8403
rect 4244 8351 4300 8383
rect 4352 8351 4408 8383
rect 4460 8351 4516 8403
rect 4595 8383 4624 8403
rect 4568 8351 4624 8383
rect 4676 8383 4681 8403
rect 4784 8383 4823 8403
rect 4676 8351 4732 8383
rect 4784 8351 4840 8383
rect 4892 8351 4948 8403
rect 5021 8383 5056 8403
rect 5163 8383 5164 8403
rect 5000 8351 5056 8383
rect 5108 8351 5164 8383
rect 5216 8383 5249 8403
rect 5216 8351 5272 8383
rect 5324 8351 5380 8403
rect 5447 8383 5533 8439
rect 5589 8413 5675 8439
rect 5731 8413 5817 8439
rect 5621 8383 5675 8413
rect 5731 8383 5785 8413
rect 5873 8383 5887 8439
rect 5432 8361 5569 8383
rect 5621 8361 5677 8383
rect 5729 8361 5785 8383
rect 5837 8361 5887 8383
rect 5432 8351 5887 8361
rect 3316 8305 5887 8351
rect 3316 8297 5569 8305
rect 5621 8297 5677 8305
rect 5729 8297 5785 8305
rect 5837 8297 5887 8305
rect 3316 8295 3403 8297
rect 3459 8295 3545 8297
rect 3601 8295 3687 8297
rect 3743 8295 3829 8297
rect 3885 8295 3971 8297
rect 4027 8295 4113 8297
rect 4169 8295 4255 8297
rect 4311 8295 4397 8297
rect 4453 8295 4539 8297
rect 4595 8295 4681 8297
rect 4737 8295 4823 8297
rect 4879 8295 4965 8297
rect 5021 8295 5107 8297
rect 5163 8295 5249 8297
rect 5305 8295 5391 8297
rect 3316 8243 3328 8295
rect 3380 8243 3403 8295
rect 3488 8243 3544 8295
rect 3601 8243 3652 8295
rect 3743 8243 3760 8295
rect 3812 8243 3829 8295
rect 3920 8243 3971 8295
rect 4028 8243 4084 8295
rect 4169 8243 4192 8295
rect 4244 8243 4255 8295
rect 4352 8243 4397 8295
rect 4460 8243 4516 8295
rect 4595 8243 4624 8295
rect 4676 8243 4681 8295
rect 4784 8243 4823 8295
rect 4892 8243 4948 8295
rect 5021 8243 5056 8295
rect 5163 8243 5164 8295
rect 5216 8243 5249 8295
rect 5324 8243 5380 8295
rect 3316 8241 3403 8243
rect 3459 8241 3545 8243
rect 3601 8241 3687 8243
rect 3743 8241 3829 8243
rect 3885 8241 3971 8243
rect 4027 8241 4113 8243
rect 4169 8241 4255 8243
rect 4311 8241 4397 8243
rect 4453 8241 4539 8243
rect 4595 8241 4681 8243
rect 4737 8241 4823 8243
rect 4879 8241 4965 8243
rect 5021 8241 5107 8243
rect 5163 8241 5249 8243
rect 5305 8241 5391 8243
rect 5447 8241 5533 8297
rect 5621 8253 5675 8297
rect 5731 8253 5785 8297
rect 5589 8241 5675 8253
rect 5731 8241 5817 8253
rect 5873 8241 5887 8297
rect 3316 8197 5887 8241
rect 3316 8187 5569 8197
rect 3316 8135 3328 8187
rect 3380 8155 3436 8187
rect 3380 8135 3403 8155
rect 3488 8135 3544 8187
rect 3596 8155 3652 8187
rect 3704 8155 3760 8187
rect 3601 8135 3652 8155
rect 3743 8135 3760 8155
rect 3812 8155 3868 8187
rect 3920 8155 3976 8187
rect 3812 8135 3829 8155
rect 3920 8135 3971 8155
rect 4028 8135 4084 8187
rect 4136 8155 4192 8187
rect 4169 8135 4192 8155
rect 4244 8155 4300 8187
rect 4352 8155 4408 8187
rect 4244 8135 4255 8155
rect 4352 8135 4397 8155
rect 4460 8135 4516 8187
rect 4568 8155 4624 8187
rect 4595 8135 4624 8155
rect 4676 8155 4732 8187
rect 4784 8155 4840 8187
rect 4676 8135 4681 8155
rect 4784 8135 4823 8155
rect 4892 8135 4948 8187
rect 5000 8155 5056 8187
rect 5108 8155 5164 8187
rect 5021 8135 5056 8155
rect 5163 8135 5164 8155
rect 5216 8155 5272 8187
rect 5216 8135 5249 8155
rect 5324 8135 5380 8187
rect 5432 8155 5569 8187
rect 5621 8155 5677 8197
rect 5729 8155 5785 8197
rect 5837 8155 5887 8197
rect 3316 8099 3403 8135
rect 3459 8099 3545 8135
rect 3601 8099 3687 8135
rect 3743 8099 3829 8135
rect 3885 8099 3971 8135
rect 4027 8099 4113 8135
rect 4169 8099 4255 8135
rect 4311 8099 4397 8135
rect 4453 8099 4539 8135
rect 4595 8099 4681 8135
rect 4737 8099 4823 8135
rect 4879 8099 4965 8135
rect 5021 8099 5107 8135
rect 5163 8099 5249 8135
rect 5305 8099 5391 8135
rect 5447 8099 5533 8155
rect 5621 8145 5675 8155
rect 5731 8145 5785 8155
rect 5589 8099 5675 8145
rect 5731 8099 5817 8145
rect 5873 8099 5887 8155
rect 3316 8089 5887 8099
rect 3316 8085 5569 8089
rect 329 8037 379 8085
rect 11 7981 379 8037
rect 11 7929 61 7981
rect 113 7929 169 7981
rect 221 7929 277 7981
rect 329 7929 379 7981
rect 5519 8037 5569 8085
rect 5621 8037 5677 8089
rect 5729 8037 5785 8089
rect 5837 8037 5887 8089
rect 5519 7981 5887 8037
rect 11 7873 379 7929
rect 11 7835 61 7873
rect 113 7835 169 7873
rect 221 7835 277 7873
rect 329 7835 379 7873
rect 11 7779 25 7835
rect 113 7821 167 7835
rect 223 7821 277 7835
rect 81 7779 167 7821
rect 223 7779 309 7821
rect 365 7779 379 7835
rect 1766 7949 4130 7961
rect 1766 7793 1778 7949
rect 4118 7793 4130 7949
rect 1766 7781 4130 7793
rect 5519 7929 5569 7981
rect 5621 7929 5677 7981
rect 5729 7929 5785 7981
rect 5837 7929 5887 7981
rect 5519 7873 5887 7929
rect 5519 7835 5569 7873
rect 5621 7835 5677 7873
rect 5729 7835 5785 7873
rect 5837 7835 5887 7873
rect 11 7765 379 7779
rect 11 7713 61 7765
rect 113 7713 169 7765
rect 221 7713 277 7765
rect 329 7713 379 7765
rect 11 7693 379 7713
rect 11 7637 25 7693
rect 81 7657 167 7693
rect 223 7657 309 7693
rect 113 7637 167 7657
rect 223 7637 277 7657
rect 365 7637 379 7693
rect 11 7605 61 7637
rect 113 7605 169 7637
rect 221 7605 277 7637
rect 329 7605 379 7637
rect 11 7551 379 7605
rect 11 7495 25 7551
rect 81 7549 167 7551
rect 223 7549 309 7551
rect 113 7497 167 7549
rect 223 7497 277 7549
rect 81 7495 167 7497
rect 223 7495 309 7497
rect 365 7495 379 7551
rect 11 7441 379 7495
rect 11 7409 61 7441
rect 113 7409 169 7441
rect 221 7409 277 7441
rect 329 7409 379 7441
rect 11 7353 25 7409
rect 113 7389 167 7409
rect 223 7389 277 7409
rect 81 7353 167 7389
rect 223 7353 309 7389
rect 365 7353 379 7409
rect 11 7333 379 7353
rect 11 7281 61 7333
rect 113 7281 169 7333
rect 221 7281 277 7333
rect 329 7281 379 7333
rect 11 7267 379 7281
rect 11 7211 25 7267
rect 81 7225 167 7267
rect 223 7225 309 7267
rect 113 7211 167 7225
rect 223 7211 277 7225
rect 365 7211 379 7267
rect 11 7173 61 7211
rect 113 7173 169 7211
rect 221 7173 277 7211
rect 329 7173 379 7211
rect 11 7125 379 7173
rect 5519 7779 5533 7835
rect 5621 7821 5675 7835
rect 5731 7821 5785 7835
rect 5589 7779 5675 7821
rect 5731 7779 5817 7821
rect 5873 7779 5887 7835
rect 5519 7765 5887 7779
rect 5519 7713 5569 7765
rect 5621 7713 5677 7765
rect 5729 7713 5785 7765
rect 5837 7713 5887 7765
rect 5519 7693 5887 7713
rect 5519 7637 5533 7693
rect 5589 7657 5675 7693
rect 5731 7657 5817 7693
rect 5621 7637 5675 7657
rect 5731 7637 5785 7657
rect 5873 7637 5887 7693
rect 5519 7605 5569 7637
rect 5621 7605 5677 7637
rect 5729 7605 5785 7637
rect 5837 7605 5887 7637
rect 5519 7551 5887 7605
rect 5519 7495 5533 7551
rect 5589 7549 5675 7551
rect 5731 7549 5817 7551
rect 5621 7497 5675 7549
rect 5731 7497 5785 7549
rect 5589 7495 5675 7497
rect 5731 7495 5817 7497
rect 5873 7495 5887 7551
rect 5519 7441 5887 7495
rect 5519 7409 5569 7441
rect 5621 7409 5677 7441
rect 5729 7409 5785 7441
rect 5837 7409 5887 7441
rect 5519 7353 5533 7409
rect 5621 7389 5675 7409
rect 5731 7389 5785 7409
rect 5589 7353 5675 7389
rect 5731 7353 5817 7389
rect 5873 7353 5887 7409
rect 5519 7333 5887 7353
rect 5519 7281 5569 7333
rect 5621 7281 5677 7333
rect 5729 7281 5785 7333
rect 5837 7281 5887 7333
rect 5519 7267 5887 7281
rect 5519 7211 5533 7267
rect 5589 7225 5675 7267
rect 5731 7225 5817 7267
rect 5621 7211 5675 7225
rect 5731 7211 5785 7225
rect 5873 7211 5887 7267
rect 5519 7173 5569 7211
rect 5621 7173 5677 7211
rect 5729 7173 5785 7211
rect 5837 7173 5887 7211
rect 11 7069 25 7125
rect 81 7117 167 7125
rect 223 7117 309 7125
rect 113 7069 167 7117
rect 223 7069 277 7117
rect 365 7069 379 7125
rect 11 7065 61 7069
rect 113 7065 169 7069
rect 221 7065 277 7069
rect 329 7065 379 7069
rect 11 7009 379 7065
rect 11 6983 61 7009
rect 113 6983 169 7009
rect 221 6983 277 7009
rect 329 6983 379 7009
rect 11 6927 25 6983
rect 113 6957 167 6983
rect 223 6957 277 6983
rect 81 6927 167 6957
rect 223 6927 309 6957
rect 365 6927 379 6983
rect 11 6901 379 6927
rect 11 6849 61 6901
rect 113 6849 169 6901
rect 221 6849 277 6901
rect 329 6849 379 6901
rect 11 6841 379 6849
rect 11 6785 25 6841
rect 81 6793 167 6841
rect 223 6793 309 6841
rect 113 6785 167 6793
rect 223 6785 277 6793
rect 365 6785 379 6841
rect 11 6741 61 6785
rect 113 6741 169 6785
rect 221 6741 277 6785
rect 329 6741 379 6785
rect 11 6699 379 6741
rect 11 6643 25 6699
rect 81 6685 167 6699
rect 223 6685 309 6699
rect 113 6643 167 6685
rect 223 6643 277 6685
rect 365 6643 379 6699
rect 11 6633 61 6643
rect 113 6633 169 6643
rect 221 6633 277 6643
rect 329 6633 379 6643
rect 11 6577 379 6633
rect 11 6557 61 6577
rect 113 6557 169 6577
rect 221 6557 277 6577
rect 329 6557 379 6577
rect 11 6501 25 6557
rect 113 6525 167 6557
rect 223 6525 277 6557
rect 81 6501 167 6525
rect 223 6501 309 6525
rect 365 6501 379 6557
rect 11 6485 379 6501
rect 949 7145 4949 7157
rect 949 6989 1778 7145
rect 4118 6989 4949 7145
rect 949 6485 4949 6989
rect 5519 7125 5887 7173
rect 5519 7069 5533 7125
rect 5589 7117 5675 7125
rect 5731 7117 5817 7125
rect 5621 7069 5675 7117
rect 5731 7069 5785 7117
rect 5873 7069 5887 7125
rect 5519 7065 5569 7069
rect 5621 7065 5677 7069
rect 5729 7065 5785 7069
rect 5837 7065 5887 7069
rect 5519 7009 5887 7065
rect 5519 6983 5569 7009
rect 5621 6983 5677 7009
rect 5729 6983 5785 7009
rect 5837 6983 5887 7009
rect 5519 6927 5533 6983
rect 5621 6957 5675 6983
rect 5731 6957 5785 6983
rect 5589 6927 5675 6957
rect 5731 6927 5817 6957
rect 5873 6927 5887 6983
rect 5519 6901 5887 6927
rect 5519 6849 5569 6901
rect 5621 6849 5677 6901
rect 5729 6849 5785 6901
rect 5837 6849 5887 6901
rect 5519 6841 5887 6849
rect 5519 6785 5533 6841
rect 5589 6793 5675 6841
rect 5731 6793 5817 6841
rect 5621 6785 5675 6793
rect 5731 6785 5785 6793
rect 5873 6785 5887 6841
rect 5519 6741 5569 6785
rect 5621 6741 5677 6785
rect 5729 6741 5785 6785
rect 5837 6741 5887 6785
rect 5519 6699 5887 6741
rect 5519 6643 5533 6699
rect 5589 6685 5675 6699
rect 5731 6685 5817 6699
rect 5621 6643 5675 6685
rect 5731 6643 5785 6685
rect 5873 6643 5887 6699
rect 5519 6633 5569 6643
rect 5621 6633 5677 6643
rect 5729 6633 5785 6643
rect 5837 6633 5887 6643
rect 5519 6577 5887 6633
rect 5519 6557 5569 6577
rect 5621 6557 5677 6577
rect 5729 6557 5785 6577
rect 5837 6557 5887 6577
rect 5519 6501 5533 6557
rect 5621 6525 5675 6557
rect 5731 6525 5785 6557
rect 5589 6501 5675 6525
rect 5731 6501 5817 6525
rect 5873 6501 5887 6557
rect 5519 6485 5887 6501
rect 548 5708 770 5750
rect 548 5688 579 5708
rect 548 5632 560 5688
rect 631 5656 687 5708
rect 739 5688 770 5708
rect 616 5632 702 5656
rect 758 5632 770 5688
rect 548 5600 770 5632
rect 548 5548 579 5600
rect 631 5548 687 5600
rect 739 5548 770 5600
rect 548 5546 770 5548
rect 548 5490 560 5546
rect 616 5492 702 5546
rect 548 5440 579 5490
rect 631 5440 687 5492
rect 758 5490 770 5546
rect 739 5440 770 5490
rect 548 5404 770 5440
rect 548 5348 560 5404
rect 616 5384 702 5404
rect 548 5332 579 5348
rect 631 5332 687 5384
rect 758 5348 770 5404
rect 739 5332 770 5348
rect 548 5276 770 5332
rect 548 5262 579 5276
rect 548 5206 560 5262
rect 631 5224 687 5276
rect 739 5262 770 5276
rect 616 5206 702 5224
rect 758 5206 770 5262
rect 548 5168 770 5206
rect 548 5120 579 5168
rect 548 5064 560 5120
rect 631 5116 687 5168
rect 739 5120 770 5168
rect 616 5064 702 5116
rect 758 5064 770 5120
rect 548 5060 770 5064
rect 548 5008 579 5060
rect 631 5008 687 5060
rect 739 5008 770 5060
rect 548 4978 770 5008
rect 548 4922 560 4978
rect 616 4952 702 4978
rect 548 4900 579 4922
rect 631 4900 687 4952
rect 758 4922 770 4978
rect 739 4900 770 4922
rect 548 4859 770 4900
rect 949 5327 1395 6485
rect 949 5171 990 5327
rect 1354 5171 1395 5327
rect 11 4624 379 4659
rect 11 4568 25 4624
rect 81 4611 167 4624
rect 223 4611 309 4624
rect 113 4568 167 4611
rect 223 4568 277 4611
rect 365 4568 379 4624
rect 11 4559 61 4568
rect 113 4559 169 4568
rect 221 4559 277 4568
rect 329 4559 379 4568
rect 11 4503 379 4559
rect 11 4482 61 4503
rect 113 4482 169 4503
rect 221 4482 277 4503
rect 329 4482 379 4503
rect 11 4426 25 4482
rect 113 4451 167 4482
rect 223 4451 277 4482
rect 81 4426 167 4451
rect 223 4426 309 4451
rect 365 4426 379 4482
rect 11 4395 379 4426
rect 11 4343 61 4395
rect 113 4343 169 4395
rect 221 4343 277 4395
rect 329 4343 379 4395
rect 11 4340 379 4343
rect 11 4284 25 4340
rect 81 4287 167 4340
rect 223 4287 309 4340
rect 113 4284 167 4287
rect 223 4284 277 4287
rect 365 4284 379 4340
rect 11 4235 61 4284
rect 113 4235 169 4284
rect 221 4235 277 4284
rect 329 4235 379 4284
rect 11 4198 379 4235
rect 11 4142 25 4198
rect 81 4179 167 4198
rect 223 4179 309 4198
rect 113 4142 167 4179
rect 223 4142 277 4179
rect 365 4142 379 4198
rect 11 4127 61 4142
rect 113 4127 169 4142
rect 221 4127 277 4142
rect 329 4127 379 4142
rect 11 4071 379 4127
rect 11 4056 61 4071
rect 113 4056 169 4071
rect 221 4056 277 4071
rect 329 4056 379 4071
rect 11 4000 25 4056
rect 113 4019 167 4056
rect 223 4019 277 4056
rect 81 4000 167 4019
rect 223 4000 309 4019
rect 365 4000 379 4056
rect 11 3963 379 4000
rect 11 3914 61 3963
rect 113 3914 169 3963
rect 221 3914 277 3963
rect 329 3914 379 3963
rect 11 3858 25 3914
rect 113 3911 167 3914
rect 223 3911 277 3914
rect 81 3858 167 3911
rect 223 3858 309 3911
rect 365 3858 379 3914
rect 11 3855 379 3858
rect 11 3803 61 3855
rect 113 3803 169 3855
rect 221 3803 277 3855
rect 329 3803 379 3855
rect 11 3772 379 3803
rect 11 3716 25 3772
rect 81 3747 167 3772
rect 223 3747 309 3772
rect 113 3716 167 3747
rect 223 3716 277 3747
rect 365 3716 379 3772
rect 11 3695 61 3716
rect 113 3695 169 3716
rect 221 3695 277 3716
rect 329 3695 379 3716
rect 11 3639 379 3695
rect 11 3630 61 3639
rect 113 3630 169 3639
rect 221 3630 277 3639
rect 329 3630 379 3639
rect 11 3574 25 3630
rect 113 3587 167 3630
rect 223 3587 277 3630
rect 81 3574 167 3587
rect 223 3574 309 3587
rect 365 3574 379 3630
rect 11 3539 379 3574
rect 949 4393 1395 5171
rect 949 4237 990 4393
rect 1354 4237 1395 4393
rect 949 3439 1395 4237
rect 1455 5717 1901 5750
rect 1455 5561 1496 5717
rect 1860 5561 1901 5717
rect 1455 5546 1901 5561
rect 1455 5490 1508 5546
rect 1564 5490 1650 5546
rect 1706 5490 1792 5546
rect 1848 5490 1901 5546
rect 1455 5404 1901 5490
rect 1455 5348 1508 5404
rect 1564 5348 1650 5404
rect 1706 5348 1792 5404
rect 1848 5348 1901 5404
rect 1455 5262 1901 5348
rect 1455 5206 1508 5262
rect 1564 5206 1650 5262
rect 1706 5206 1792 5262
rect 1848 5206 1901 5262
rect 1455 5120 1901 5206
rect 1455 5064 1508 5120
rect 1564 5064 1650 5120
rect 1706 5064 1792 5120
rect 1848 5064 1901 5120
rect 1455 4978 1901 5064
rect 1455 4922 1508 4978
rect 1564 4922 1650 4978
rect 1706 4922 1792 4978
rect 1848 4922 1901 4978
rect 1455 4912 1901 4922
rect 1455 4652 1496 4912
rect 1860 4652 1901 4912
rect 1455 4003 1901 4652
rect 1455 3847 1496 4003
rect 1860 3847 1901 4003
rect 1455 3814 1901 3847
rect 1961 5327 2407 6485
rect 1961 5171 2002 5327
rect 2366 5171 2407 5327
rect 1961 4393 2407 5171
rect 1961 4237 2002 4393
rect 2366 4237 2407 4393
rect 1961 3439 2407 4237
rect 2467 5717 2913 5750
rect 2467 5561 2508 5717
rect 2872 5561 2913 5717
rect 2467 5546 2913 5561
rect 2467 5490 2520 5546
rect 2576 5490 2662 5546
rect 2718 5490 2804 5546
rect 2860 5490 2913 5546
rect 2467 5404 2913 5490
rect 2467 5348 2520 5404
rect 2576 5348 2662 5404
rect 2718 5348 2804 5404
rect 2860 5348 2913 5404
rect 2467 5262 2913 5348
rect 2467 5206 2520 5262
rect 2576 5206 2662 5262
rect 2718 5206 2804 5262
rect 2860 5206 2913 5262
rect 2467 5120 2913 5206
rect 2467 5064 2520 5120
rect 2576 5064 2662 5120
rect 2718 5064 2804 5120
rect 2860 5064 2913 5120
rect 2467 4978 2913 5064
rect 2467 4922 2520 4978
rect 2576 4922 2662 4978
rect 2718 4922 2804 4978
rect 2860 4922 2913 4978
rect 2467 4912 2913 4922
rect 2467 4652 2508 4912
rect 2872 4652 2913 4912
rect 2467 4003 2913 4652
rect 2467 3847 2508 4003
rect 2872 3847 2913 4003
rect 2467 3814 2913 3847
rect 2985 5717 3431 5750
rect 2985 5561 3026 5717
rect 3390 5561 3431 5717
rect 2985 5546 3431 5561
rect 2985 5490 3038 5546
rect 3094 5490 3180 5546
rect 3236 5490 3322 5546
rect 3378 5490 3431 5546
rect 2985 5404 3431 5490
rect 2985 5348 3038 5404
rect 3094 5348 3180 5404
rect 3236 5348 3322 5404
rect 3378 5348 3431 5404
rect 2985 5262 3431 5348
rect 2985 5206 3038 5262
rect 3094 5206 3180 5262
rect 3236 5206 3322 5262
rect 3378 5206 3431 5262
rect 2985 5120 3431 5206
rect 2985 5064 3038 5120
rect 3094 5064 3180 5120
rect 3236 5064 3322 5120
rect 3378 5064 3431 5120
rect 2985 4978 3431 5064
rect 2985 4922 3038 4978
rect 3094 4922 3180 4978
rect 3236 4922 3322 4978
rect 3378 4922 3431 4978
rect 2985 4912 3431 4922
rect 2985 4652 3026 4912
rect 3390 4652 3431 4912
rect 2985 4003 3431 4652
rect 2985 3847 3026 4003
rect 3390 3847 3431 4003
rect 2985 3814 3431 3847
rect 3491 5327 3937 6485
rect 3491 5171 3532 5327
rect 3896 5171 3937 5327
rect 3491 4393 3937 5171
rect 3491 4237 3532 4393
rect 3896 4237 3937 4393
rect 3491 3439 3937 4237
rect 3997 5717 4443 5750
rect 3997 5561 4038 5717
rect 4402 5561 4443 5717
rect 3997 5546 4443 5561
rect 3997 5490 4050 5546
rect 4106 5490 4192 5546
rect 4248 5490 4334 5546
rect 4390 5490 4443 5546
rect 3997 5404 4443 5490
rect 3997 5348 4050 5404
rect 4106 5348 4192 5404
rect 4248 5348 4334 5404
rect 4390 5348 4443 5404
rect 3997 5262 4443 5348
rect 3997 5206 4050 5262
rect 4106 5206 4192 5262
rect 4248 5206 4334 5262
rect 4390 5206 4443 5262
rect 3997 5120 4443 5206
rect 3997 5064 4050 5120
rect 4106 5064 4192 5120
rect 4248 5064 4334 5120
rect 4390 5064 4443 5120
rect 3997 4978 4443 5064
rect 3997 4922 4050 4978
rect 4106 4922 4192 4978
rect 4248 4922 4334 4978
rect 4390 4922 4443 4978
rect 3997 4912 4443 4922
rect 3997 4652 4038 4912
rect 4402 4652 4443 4912
rect 3997 4003 4443 4652
rect 3997 3847 4038 4003
rect 4402 3847 4443 4003
rect 3997 3814 4443 3847
rect 4503 5327 4949 6485
rect 4503 5171 4544 5327
rect 4908 5171 4949 5327
rect 4503 4393 4949 5171
rect 5128 5708 5350 5750
rect 5128 5688 5159 5708
rect 5128 5632 5140 5688
rect 5211 5656 5267 5708
rect 5319 5688 5350 5708
rect 5196 5632 5282 5656
rect 5338 5632 5350 5688
rect 5128 5600 5350 5632
rect 5128 5548 5159 5600
rect 5211 5548 5267 5600
rect 5319 5548 5350 5600
rect 5128 5546 5350 5548
rect 5128 5490 5140 5546
rect 5196 5492 5282 5546
rect 5128 5440 5159 5490
rect 5211 5440 5267 5492
rect 5338 5490 5350 5546
rect 5319 5440 5350 5490
rect 5128 5404 5350 5440
rect 5128 5348 5140 5404
rect 5196 5384 5282 5404
rect 5128 5332 5159 5348
rect 5211 5332 5267 5384
rect 5338 5348 5350 5404
rect 5319 5332 5350 5348
rect 5128 5276 5350 5332
rect 5128 5262 5159 5276
rect 5128 5206 5140 5262
rect 5211 5224 5267 5276
rect 5319 5262 5350 5276
rect 5196 5206 5282 5224
rect 5338 5206 5350 5262
rect 5128 5168 5350 5206
rect 5128 5120 5159 5168
rect 5128 5064 5140 5120
rect 5211 5116 5267 5168
rect 5319 5120 5350 5168
rect 5196 5064 5282 5116
rect 5338 5064 5350 5120
rect 5128 5060 5350 5064
rect 5128 5008 5159 5060
rect 5211 5008 5267 5060
rect 5319 5008 5350 5060
rect 5128 4978 5350 5008
rect 5128 4922 5140 4978
rect 5196 4952 5282 4978
rect 5128 4900 5159 4922
rect 5211 4900 5267 4952
rect 5338 4922 5350 4978
rect 5319 4900 5350 4922
rect 5128 4859 5350 4900
rect 4503 4237 4544 4393
rect 4908 4237 4949 4393
rect 4503 3439 4949 4237
rect -205 2939 4949 3439
rect 5519 4633 5887 4659
rect 5519 4626 5569 4633
rect 5621 4626 5677 4633
rect 5729 4626 5785 4633
rect 5837 4626 5887 4633
rect 5519 4570 5533 4626
rect 5621 4581 5675 4626
rect 5731 4581 5785 4626
rect 5589 4570 5675 4581
rect 5731 4570 5817 4581
rect 5873 4570 5887 4626
rect 5519 4525 5887 4570
rect 5519 4484 5569 4525
rect 5621 4484 5677 4525
rect 5729 4484 5785 4525
rect 5837 4484 5887 4525
rect 5519 4428 5533 4484
rect 5621 4473 5675 4484
rect 5731 4473 5785 4484
rect 5589 4428 5675 4473
rect 5731 4428 5817 4473
rect 5873 4428 5887 4484
rect 5519 4417 5887 4428
rect 5519 4365 5569 4417
rect 5621 4365 5677 4417
rect 5729 4365 5785 4417
rect 5837 4365 5887 4417
rect 5519 4342 5887 4365
rect 5519 4286 5533 4342
rect 5589 4309 5675 4342
rect 5731 4309 5817 4342
rect 5621 4286 5675 4309
rect 5731 4286 5785 4309
rect 5873 4286 5887 4342
rect 5519 4257 5569 4286
rect 5621 4257 5677 4286
rect 5729 4257 5785 4286
rect 5837 4257 5887 4286
rect 5519 4201 5887 4257
rect 5519 4200 5569 4201
rect 5621 4200 5677 4201
rect 5729 4200 5785 4201
rect 5837 4200 5887 4201
rect 5519 4144 5533 4200
rect 5621 4149 5675 4200
rect 5731 4149 5785 4200
rect 5589 4144 5675 4149
rect 5731 4144 5817 4149
rect 5873 4144 5887 4200
rect 5519 4093 5887 4144
rect 5519 4058 5569 4093
rect 5621 4058 5677 4093
rect 5729 4058 5785 4093
rect 5837 4058 5887 4093
rect 5519 4002 5533 4058
rect 5621 4041 5675 4058
rect 5731 4041 5785 4058
rect 5589 4002 5675 4041
rect 5731 4002 5817 4041
rect 5873 4002 5887 4058
rect 5519 3985 5887 4002
rect 5519 3933 5569 3985
rect 5621 3933 5677 3985
rect 5729 3933 5785 3985
rect 5837 3933 5887 3985
rect 5519 3916 5887 3933
rect 5519 3860 5533 3916
rect 5589 3877 5675 3916
rect 5731 3877 5817 3916
rect 5621 3860 5675 3877
rect 5731 3860 5785 3877
rect 5873 3860 5887 3916
rect 5519 3825 5569 3860
rect 5621 3825 5677 3860
rect 5729 3825 5785 3860
rect 5837 3825 5887 3860
rect 5519 3774 5887 3825
rect 5519 3718 5533 3774
rect 5589 3769 5675 3774
rect 5731 3769 5817 3774
rect 5621 3718 5675 3769
rect 5731 3718 5785 3769
rect 5873 3718 5887 3774
rect 5519 3717 5569 3718
rect 5621 3717 5677 3718
rect 5729 3717 5785 3718
rect 5837 3717 5887 3718
rect 5519 3661 5887 3717
rect 5519 3632 5569 3661
rect 5621 3632 5677 3661
rect 5729 3632 5785 3661
rect 5837 3632 5887 3661
rect 5519 3576 5533 3632
rect 5621 3609 5675 3632
rect 5731 3609 5785 3632
rect 5589 3576 5675 3609
rect 5731 3576 5817 3609
rect 5873 3576 5887 3632
rect 5519 3553 5887 3576
rect 5519 3501 5569 3553
rect 5621 3501 5677 3553
rect 5729 3501 5785 3553
rect 5837 3501 5887 3553
rect 5519 3490 5887 3501
rect 5519 3434 5533 3490
rect 5589 3445 5675 3490
rect 5731 3445 5817 3490
rect 5621 3434 5675 3445
rect 5731 3434 5785 3445
rect 5873 3434 5887 3490
rect 5519 3393 5569 3434
rect 5621 3393 5677 3434
rect 5729 3393 5785 3434
rect 5837 3393 5887 3434
rect 5519 3348 5887 3393
rect 5519 3292 5533 3348
rect 5589 3337 5675 3348
rect 5731 3337 5817 3348
rect 5621 3292 5675 3337
rect 5731 3292 5785 3337
rect 5873 3292 5887 3348
rect 5519 3285 5569 3292
rect 5621 3285 5677 3292
rect 5729 3285 5785 3292
rect 5837 3285 5887 3292
rect 5519 3259 5887 3285
rect 11 2821 379 2839
rect 11 2779 61 2821
rect 113 2779 169 2821
rect 221 2779 277 2821
rect 329 2779 379 2821
rect 11 2723 25 2779
rect 113 2769 167 2779
rect 223 2769 277 2779
rect 81 2723 167 2769
rect 223 2723 309 2769
rect 365 2723 379 2779
rect 11 2713 379 2723
rect 11 2661 61 2713
rect 113 2661 169 2713
rect 221 2661 277 2713
rect 329 2661 379 2713
rect 11 2637 379 2661
rect 11 2581 25 2637
rect 81 2605 167 2637
rect 223 2605 309 2637
rect 113 2581 167 2605
rect 223 2581 277 2605
rect 365 2581 379 2637
rect 11 2553 61 2581
rect 113 2553 169 2581
rect 221 2553 277 2581
rect 329 2553 379 2581
rect 11 2497 379 2553
rect 11 2495 61 2497
rect 113 2495 169 2497
rect 221 2495 277 2497
rect 329 2495 379 2497
rect 11 2439 25 2495
rect 113 2445 167 2495
rect 223 2445 277 2495
rect 81 2439 167 2445
rect 223 2439 309 2445
rect 365 2439 379 2495
rect 11 2389 379 2439
rect 11 2353 61 2389
rect 113 2353 169 2389
rect 221 2353 277 2389
rect 329 2353 379 2389
rect 11 2297 25 2353
rect 113 2337 167 2353
rect 223 2337 277 2353
rect 81 2297 167 2337
rect 223 2297 309 2337
rect 365 2297 379 2353
rect 11 2281 379 2297
rect 11 2229 61 2281
rect 113 2229 169 2281
rect 221 2229 277 2281
rect 329 2229 379 2281
rect 11 2211 379 2229
rect 11 2155 25 2211
rect 81 2173 167 2211
rect 223 2173 309 2211
rect 113 2155 167 2173
rect 223 2155 277 2173
rect 365 2155 379 2211
rect 11 2121 61 2155
rect 113 2121 169 2155
rect 221 2121 277 2155
rect 329 2121 379 2155
rect 11 2069 379 2121
rect 11 2013 25 2069
rect 81 2065 167 2069
rect 223 2065 309 2069
rect 113 2013 167 2065
rect 223 2013 277 2065
rect 365 2013 379 2069
rect 11 1957 379 2013
rect 11 1927 61 1957
rect 113 1927 169 1957
rect 221 1927 277 1957
rect 329 1927 379 1957
rect 11 1871 25 1927
rect 113 1905 167 1927
rect 223 1905 277 1927
rect 81 1871 167 1905
rect 223 1871 309 1905
rect 365 1871 379 1927
rect 11 1849 379 1871
rect 11 1797 61 1849
rect 113 1797 169 1849
rect 221 1797 277 1849
rect 329 1797 379 1849
rect 11 1785 379 1797
rect 11 1729 25 1785
rect 81 1741 167 1785
rect 223 1741 309 1785
rect 113 1729 167 1741
rect 223 1729 277 1741
rect 365 1729 379 1785
rect 11 1689 61 1729
rect 113 1689 169 1729
rect 221 1689 277 1729
rect 329 1689 379 1729
rect 11 1659 379 1689
rect 949 2090 1395 2939
rect 949 1934 990 2090
rect 1354 1934 1395 2090
rect 548 1418 770 1428
rect 548 1362 560 1418
rect 616 1416 702 1418
rect 631 1364 687 1416
rect 616 1362 702 1364
rect 758 1362 770 1418
rect 548 1308 770 1362
rect 548 1276 579 1308
rect 548 1220 560 1276
rect 631 1256 687 1308
rect 739 1276 770 1308
rect 616 1220 702 1256
rect 758 1220 770 1276
rect 548 1200 770 1220
rect 548 1148 579 1200
rect 631 1148 687 1200
rect 739 1148 770 1200
rect 548 1134 770 1148
rect 548 1078 560 1134
rect 616 1092 702 1134
rect 548 1040 579 1078
rect 631 1040 687 1092
rect 758 1078 770 1134
rect 739 1040 770 1078
rect 548 992 770 1040
rect 548 936 560 992
rect 616 984 702 992
rect 548 932 579 936
rect 631 932 687 984
rect 758 936 770 992
rect 949 1156 1395 1934
rect 949 1000 990 1156
rect 1354 1000 1395 1156
rect 949 978 1395 1000
rect 1455 2480 1901 2513
rect 1455 2324 1496 2480
rect 1860 2324 1901 2480
rect 1455 1675 1901 2324
rect 1455 1415 1496 1675
rect 1860 1415 1901 1675
rect 1455 1362 1508 1415
rect 1564 1362 1650 1415
rect 1706 1362 1792 1415
rect 1848 1362 1901 1415
rect 1455 1276 1901 1362
rect 1455 1220 1508 1276
rect 1564 1220 1650 1276
rect 1706 1220 1792 1276
rect 1848 1220 1901 1276
rect 1455 1134 1901 1220
rect 1455 1078 1508 1134
rect 1564 1078 1650 1134
rect 1706 1078 1792 1134
rect 1848 1078 1901 1134
rect 1455 992 1901 1078
rect 739 932 770 936
rect 548 876 770 932
rect 548 824 579 876
rect 631 824 687 876
rect 739 824 770 876
rect 548 797 770 824
rect 1455 936 1508 992
rect 1564 936 1650 992
rect 1706 936 1792 992
rect 1848 936 1901 992
rect 1961 2090 2407 2939
rect 1961 1934 2002 2090
rect 2366 1934 2407 2090
rect 1961 1156 2407 1934
rect 1961 1000 2002 1156
rect 2366 1000 2407 1156
rect 1961 978 2407 1000
rect 2514 2480 2754 2513
rect 2514 2324 2556 2480
rect 2712 2324 2754 2480
rect 2514 1675 2754 2324
rect 2514 1418 2554 1675
rect 2710 1418 2754 1675
rect 2514 1362 2535 1418
rect 2591 1362 2677 1415
rect 2733 1362 2754 1418
rect 2514 1276 2754 1362
rect 2514 1220 2535 1276
rect 2591 1220 2677 1276
rect 2733 1220 2754 1276
rect 2514 1134 2754 1220
rect 2514 1078 2535 1134
rect 2591 1078 2677 1134
rect 2733 1078 2754 1134
rect 2514 992 2754 1078
rect 1455 797 1901 936
rect 2514 936 2535 992
rect 2591 936 2677 992
rect 2733 936 2754 992
rect 2514 797 2754 936
rect 3145 2480 3385 2513
rect 3145 2324 3187 2480
rect 3343 2324 3385 2480
rect 3145 1675 3385 2324
rect 3145 1418 3185 1675
rect 3341 1418 3385 1675
rect 3145 1362 3166 1418
rect 3222 1362 3308 1415
rect 3364 1362 3385 1418
rect 3145 1276 3385 1362
rect 3145 1220 3166 1276
rect 3222 1220 3308 1276
rect 3364 1220 3385 1276
rect 3145 1134 3385 1220
rect 3145 1078 3166 1134
rect 3222 1078 3308 1134
rect 3364 1078 3385 1134
rect 3145 992 3385 1078
rect 3145 936 3166 992
rect 3222 936 3308 992
rect 3364 936 3385 992
rect 3491 2090 3937 2939
rect 3491 1934 3532 2090
rect 3896 1934 3937 2090
rect 3491 1156 3937 1934
rect 3491 1000 3532 1156
rect 3896 1000 3937 1156
rect 3491 978 3937 1000
rect 3997 2480 4443 2513
rect 3997 2324 4038 2480
rect 4402 2324 4443 2480
rect 3997 1675 4443 2324
rect 3997 1415 4038 1675
rect 4402 1415 4443 1675
rect 3997 1362 4050 1415
rect 4106 1362 4192 1415
rect 4248 1362 4334 1415
rect 4390 1362 4443 1415
rect 3997 1276 4443 1362
rect 3997 1220 4050 1276
rect 4106 1220 4192 1276
rect 4248 1220 4334 1276
rect 4390 1220 4443 1276
rect 3997 1134 4443 1220
rect 3997 1078 4050 1134
rect 4106 1078 4192 1134
rect 4248 1078 4334 1134
rect 4390 1078 4443 1134
rect 3997 992 4443 1078
rect 3145 797 3385 936
rect 3997 936 4050 992
rect 4106 936 4192 992
rect 4248 936 4334 992
rect 4390 936 4443 992
rect 4503 2090 4949 2939
rect 4503 1934 4544 2090
rect 4908 1934 4949 2090
rect 4503 1156 4949 1934
rect 5519 3033 5887 3059
rect 5519 2977 5533 3033
rect 5621 2981 5675 3033
rect 5731 2981 5785 3033
rect 5589 2977 5675 2981
rect 5731 2977 5817 2981
rect 5873 2977 5887 3033
rect 5519 2925 5887 2977
rect 5519 2891 5569 2925
rect 5621 2891 5677 2925
rect 5729 2891 5785 2925
rect 5837 2891 5887 2925
rect 5519 2835 5533 2891
rect 5621 2873 5675 2891
rect 5731 2873 5785 2891
rect 5589 2835 5675 2873
rect 5731 2835 5817 2873
rect 5873 2835 5887 2891
rect 5519 2817 5887 2835
rect 5519 2765 5569 2817
rect 5621 2765 5677 2817
rect 5729 2765 5785 2817
rect 5837 2765 5887 2817
rect 5519 2749 5887 2765
rect 5519 2693 5533 2749
rect 5589 2709 5675 2749
rect 5731 2709 5817 2749
rect 5621 2693 5675 2709
rect 5731 2693 5785 2709
rect 5873 2693 5887 2749
rect 5519 2657 5569 2693
rect 5621 2657 5677 2693
rect 5729 2657 5785 2693
rect 5837 2657 5887 2693
rect 5519 2607 5887 2657
rect 5519 2551 5533 2607
rect 5589 2601 5675 2607
rect 5731 2601 5817 2607
rect 5621 2551 5675 2601
rect 5731 2551 5785 2601
rect 5873 2551 5887 2607
rect 5519 2549 5569 2551
rect 5621 2549 5677 2551
rect 5729 2549 5785 2551
rect 5837 2549 5887 2551
rect 5519 2493 5887 2549
rect 5519 2465 5569 2493
rect 5621 2465 5677 2493
rect 5729 2465 5785 2493
rect 5837 2465 5887 2493
rect 5519 2409 5533 2465
rect 5621 2441 5675 2465
rect 5731 2441 5785 2465
rect 5589 2409 5675 2441
rect 5731 2409 5817 2441
rect 5873 2409 5887 2465
rect 5519 2385 5887 2409
rect 5519 2333 5569 2385
rect 5621 2333 5677 2385
rect 5729 2333 5785 2385
rect 5837 2333 5887 2385
rect 5519 2323 5887 2333
rect 5519 2267 5533 2323
rect 5589 2277 5675 2323
rect 5731 2277 5817 2323
rect 5621 2267 5675 2277
rect 5731 2267 5785 2277
rect 5873 2267 5887 2323
rect 5519 2225 5569 2267
rect 5621 2225 5677 2267
rect 5729 2225 5785 2267
rect 5837 2225 5887 2267
rect 5519 2181 5887 2225
rect 5519 2125 5533 2181
rect 5589 2169 5675 2181
rect 5731 2169 5817 2181
rect 5621 2125 5675 2169
rect 5731 2125 5785 2169
rect 5873 2125 5887 2181
rect 5519 2117 5569 2125
rect 5621 2117 5677 2125
rect 5729 2117 5785 2125
rect 5837 2117 5887 2125
rect 5519 2061 5887 2117
rect 5519 2039 5569 2061
rect 5621 2039 5677 2061
rect 5729 2039 5785 2061
rect 5837 2039 5887 2061
rect 5519 1983 5533 2039
rect 5621 2009 5675 2039
rect 5731 2009 5785 2039
rect 5589 1983 5675 2009
rect 5731 1983 5817 2009
rect 5873 1983 5887 2039
rect 5519 1953 5887 1983
rect 5519 1901 5569 1953
rect 5621 1901 5677 1953
rect 5729 1901 5785 1953
rect 5837 1901 5887 1953
rect 5519 1897 5887 1901
rect 5519 1841 5533 1897
rect 5589 1845 5675 1897
rect 5731 1845 5817 1897
rect 5621 1841 5675 1845
rect 5731 1841 5785 1845
rect 5873 1841 5887 1897
rect 5519 1793 5569 1841
rect 5621 1793 5677 1841
rect 5729 1793 5785 1841
rect 5837 1793 5887 1841
rect 5519 1755 5887 1793
rect 5519 1699 5533 1755
rect 5589 1737 5675 1755
rect 5731 1737 5817 1755
rect 5621 1699 5675 1737
rect 5731 1699 5785 1737
rect 5873 1699 5887 1755
rect 5519 1685 5569 1699
rect 5621 1685 5677 1699
rect 5729 1685 5785 1699
rect 5837 1685 5887 1699
rect 5519 1659 5887 1685
rect 4503 1000 4544 1156
rect 4908 1000 4949 1156
rect 4503 978 4949 1000
rect 5130 1418 5348 1428
rect 5130 1362 5140 1418
rect 5196 1416 5282 1418
rect 5211 1364 5267 1416
rect 5196 1362 5282 1364
rect 5338 1362 5348 1418
rect 5130 1308 5348 1362
rect 5130 1276 5159 1308
rect 5130 1220 5140 1276
rect 5211 1256 5267 1308
rect 5319 1276 5348 1308
rect 5196 1220 5282 1256
rect 5338 1220 5348 1276
rect 5130 1200 5348 1220
rect 5130 1148 5159 1200
rect 5211 1148 5267 1200
rect 5319 1148 5348 1200
rect 5130 1134 5348 1148
rect 5130 1078 5140 1134
rect 5196 1092 5282 1134
rect 5130 1040 5159 1078
rect 5211 1040 5267 1092
rect 5338 1078 5348 1134
rect 5319 1040 5348 1078
rect 5130 992 5348 1040
rect 3997 797 4443 936
rect 5130 936 5140 992
rect 5196 984 5282 992
rect 5130 932 5159 936
rect 5211 932 5267 984
rect 5338 936 5348 992
rect 5319 932 5348 936
rect 5130 876 5348 932
rect 5130 824 5159 876
rect 5211 824 5267 876
rect 5319 824 5348 876
rect 5130 797 5348 824
rect 548 787 2774 797
rect 548 731 578 787
rect 634 768 720 787
rect 776 768 862 787
rect 918 768 1004 787
rect 1060 768 1146 787
rect 1202 768 1288 787
rect 1344 768 1430 787
rect 1486 768 1572 787
rect 1628 768 1714 787
rect 1770 768 1856 787
rect 1912 768 1998 787
rect 2054 768 2140 787
rect 2196 768 2282 787
rect 2338 768 2424 787
rect 2480 768 2566 787
rect 2622 768 2708 787
rect 634 731 687 768
rect 776 731 817 768
rect 918 731 925 768
rect 548 716 579 731
rect 631 716 687 731
rect 739 716 817 731
rect 869 716 925 731
rect 977 731 1004 768
rect 977 716 1033 731
rect 1085 716 1141 768
rect 1202 731 1249 768
rect 1344 731 1357 768
rect 1193 716 1249 731
rect 1301 716 1357 731
rect 1409 731 1430 768
rect 1517 731 1572 768
rect 1628 731 1681 768
rect 1770 731 1789 768
rect 1409 716 1465 731
rect 1517 716 1573 731
rect 1625 716 1681 731
rect 1733 716 1789 731
rect 1841 731 1856 768
rect 1949 731 1998 768
rect 1841 716 1897 731
rect 1949 716 2005 731
rect 2057 716 2113 768
rect 2196 731 2221 768
rect 2165 716 2221 731
rect 2273 731 2282 768
rect 2381 731 2424 768
rect 2273 716 2329 731
rect 2381 716 2437 731
rect 2489 716 2545 768
rect 2622 731 2653 768
rect 2597 716 2653 731
rect 2705 731 2708 768
rect 2764 731 2774 787
rect 2705 716 2774 731
rect 548 660 2774 716
rect 548 645 579 660
rect 631 645 687 660
rect 739 645 817 660
rect 869 645 925 660
rect 548 589 578 645
rect 634 608 687 645
rect 776 608 817 645
rect 918 608 925 645
rect 977 645 1033 660
rect 977 608 1004 645
rect 1085 608 1141 660
rect 1193 645 1249 660
rect 1301 645 1357 660
rect 1202 608 1249 645
rect 1344 608 1357 645
rect 1409 645 1465 660
rect 1517 645 1573 660
rect 1625 645 1681 660
rect 1733 645 1789 660
rect 1409 608 1430 645
rect 1517 608 1572 645
rect 1628 608 1681 645
rect 1770 608 1789 645
rect 1841 645 1897 660
rect 1949 645 2005 660
rect 1841 608 1856 645
rect 1949 608 1998 645
rect 2057 608 2113 660
rect 2165 645 2221 660
rect 2196 608 2221 645
rect 2273 645 2329 660
rect 2381 645 2437 660
rect 2273 608 2282 645
rect 2381 608 2424 645
rect 2489 608 2545 660
rect 2597 645 2653 660
rect 2622 608 2653 645
rect 2705 645 2774 660
rect 2705 608 2708 645
rect 634 589 720 608
rect 776 589 862 608
rect 918 589 1004 608
rect 1060 589 1146 608
rect 1202 589 1288 608
rect 1344 589 1430 608
rect 1486 589 1572 608
rect 1628 589 1714 608
rect 1770 589 1856 608
rect 1912 589 1998 608
rect 2054 589 2140 608
rect 2196 589 2282 608
rect 2338 589 2424 608
rect 2480 589 2566 608
rect 2622 589 2708 608
rect 2764 589 2774 645
rect 548 579 2774 589
rect 3124 787 5348 797
rect 3124 731 3134 787
rect 3190 768 3276 787
rect 3332 768 3418 787
rect 3474 768 3560 787
rect 3616 768 3702 787
rect 3758 768 3844 787
rect 3900 768 3986 787
rect 4042 768 4128 787
rect 4184 768 4270 787
rect 4326 768 4412 787
rect 4468 768 4554 787
rect 4610 768 4696 787
rect 4752 768 4838 787
rect 4894 768 4980 787
rect 5036 768 5122 787
rect 5178 768 5264 787
rect 3190 731 3193 768
rect 3124 716 3193 731
rect 3245 731 3276 768
rect 3245 716 3301 731
rect 3353 716 3409 768
rect 3474 731 3517 768
rect 3616 731 3625 768
rect 3461 716 3517 731
rect 3569 716 3625 731
rect 3677 731 3702 768
rect 3677 716 3733 731
rect 3785 716 3841 768
rect 3900 731 3949 768
rect 4042 731 4057 768
rect 3893 716 3949 731
rect 4001 716 4057 731
rect 4109 731 4128 768
rect 4217 731 4270 768
rect 4326 731 4381 768
rect 4468 731 4489 768
rect 4109 716 4165 731
rect 4217 716 4273 731
rect 4325 716 4381 731
rect 4433 716 4489 731
rect 4541 731 4554 768
rect 4649 731 4696 768
rect 4541 716 4597 731
rect 4649 716 4705 731
rect 4757 716 4813 768
rect 4894 731 4921 768
rect 4865 716 4921 731
rect 4973 731 4980 768
rect 5081 731 5122 768
rect 5211 731 5264 768
rect 5320 731 5348 787
rect 4973 716 5029 731
rect 5081 716 5159 731
rect 5211 716 5267 731
rect 5319 716 5348 731
rect 3124 660 5348 716
rect 3124 645 3193 660
rect 3124 589 3134 645
rect 3190 608 3193 645
rect 3245 645 3301 660
rect 3245 608 3276 645
rect 3353 608 3409 660
rect 3461 645 3517 660
rect 3569 645 3625 660
rect 3474 608 3517 645
rect 3616 608 3625 645
rect 3677 645 3733 660
rect 3677 608 3702 645
rect 3785 608 3841 660
rect 3893 645 3949 660
rect 4001 645 4057 660
rect 3900 608 3949 645
rect 4042 608 4057 645
rect 4109 645 4165 660
rect 4217 645 4273 660
rect 4325 645 4381 660
rect 4433 645 4489 660
rect 4109 608 4128 645
rect 4217 608 4270 645
rect 4326 608 4381 645
rect 4468 608 4489 645
rect 4541 645 4597 660
rect 4649 645 4705 660
rect 4541 608 4554 645
rect 4649 608 4696 645
rect 4757 608 4813 660
rect 4865 645 4921 660
rect 4894 608 4921 645
rect 4973 645 5029 660
rect 5081 645 5159 660
rect 5211 645 5267 660
rect 5319 645 5348 660
rect 4973 608 4980 645
rect 5081 608 5122 645
rect 5211 608 5264 645
rect 3190 589 3276 608
rect 3332 589 3418 608
rect 3474 589 3560 608
rect 3616 589 3702 608
rect 3758 589 3844 608
rect 3900 589 3986 608
rect 4042 589 4128 608
rect 4184 589 4270 608
rect 4326 589 4412 608
rect 4468 589 4554 608
rect 4610 589 4696 608
rect 4752 589 4838 608
rect 4894 589 4980 608
rect 5036 589 5122 608
rect 5178 589 5264 608
rect 5320 589 5348 645
rect 3124 579 5348 589
<< via2 >>
rect 25 8413 81 8439
rect 167 8413 223 8439
rect 309 8413 365 8439
rect 25 8383 61 8413
rect 61 8383 81 8413
rect 167 8383 169 8413
rect 169 8383 221 8413
rect 221 8383 223 8413
rect 309 8383 329 8413
rect 329 8383 365 8413
rect 451 8403 507 8439
rect 593 8403 649 8439
rect 735 8403 791 8439
rect 877 8403 933 8439
rect 1019 8403 1075 8439
rect 1161 8403 1217 8439
rect 1303 8403 1359 8439
rect 1445 8403 1501 8439
rect 1587 8403 1643 8439
rect 1729 8403 1785 8439
rect 1871 8403 1927 8439
rect 2013 8403 2069 8439
rect 2155 8403 2211 8439
rect 2297 8403 2353 8439
rect 2439 8403 2495 8439
rect 451 8383 466 8403
rect 466 8383 507 8403
rect 593 8383 626 8403
rect 626 8383 649 8403
rect 735 8383 790 8403
rect 790 8383 791 8403
rect 877 8383 898 8403
rect 898 8383 933 8403
rect 1019 8383 1058 8403
rect 1058 8383 1075 8403
rect 1161 8383 1166 8403
rect 1166 8383 1217 8403
rect 1303 8383 1330 8403
rect 1330 8383 1359 8403
rect 1445 8383 1490 8403
rect 1490 8383 1501 8403
rect 1587 8383 1598 8403
rect 1598 8383 1643 8403
rect 1729 8383 1762 8403
rect 1762 8383 1785 8403
rect 1871 8383 1922 8403
rect 1922 8383 1927 8403
rect 2013 8383 2030 8403
rect 2030 8383 2069 8403
rect 2155 8383 2194 8403
rect 2194 8383 2211 8403
rect 2297 8383 2302 8403
rect 2302 8383 2353 8403
rect 2439 8383 2462 8403
rect 2462 8383 2495 8403
rect 25 8253 61 8297
rect 61 8253 81 8297
rect 167 8253 169 8297
rect 169 8253 221 8297
rect 221 8253 223 8297
rect 309 8253 329 8297
rect 329 8253 365 8297
rect 25 8241 81 8253
rect 167 8241 223 8253
rect 309 8241 365 8253
rect 451 8295 507 8297
rect 593 8295 649 8297
rect 735 8295 791 8297
rect 877 8295 933 8297
rect 1019 8295 1075 8297
rect 1161 8295 1217 8297
rect 1303 8295 1359 8297
rect 1445 8295 1501 8297
rect 1587 8295 1643 8297
rect 1729 8295 1785 8297
rect 1871 8295 1927 8297
rect 2013 8295 2069 8297
rect 2155 8295 2211 8297
rect 2297 8295 2353 8297
rect 2439 8295 2495 8297
rect 451 8243 466 8295
rect 466 8243 507 8295
rect 593 8243 626 8295
rect 626 8243 649 8295
rect 735 8243 790 8295
rect 790 8243 791 8295
rect 877 8243 898 8295
rect 898 8243 933 8295
rect 1019 8243 1058 8295
rect 1058 8243 1075 8295
rect 1161 8243 1166 8295
rect 1166 8243 1217 8295
rect 1303 8243 1330 8295
rect 1330 8243 1359 8295
rect 1445 8243 1490 8295
rect 1490 8243 1501 8295
rect 1587 8243 1598 8295
rect 1598 8243 1643 8295
rect 1729 8243 1762 8295
rect 1762 8243 1785 8295
rect 1871 8243 1922 8295
rect 1922 8243 1927 8295
rect 2013 8243 2030 8295
rect 2030 8243 2069 8295
rect 2155 8243 2194 8295
rect 2194 8243 2211 8295
rect 2297 8243 2302 8295
rect 2302 8243 2353 8295
rect 2439 8243 2462 8295
rect 2462 8243 2495 8295
rect 451 8241 507 8243
rect 593 8241 649 8243
rect 735 8241 791 8243
rect 877 8241 933 8243
rect 1019 8241 1075 8243
rect 1161 8241 1217 8243
rect 1303 8241 1359 8243
rect 1445 8241 1501 8243
rect 1587 8241 1643 8243
rect 1729 8241 1785 8243
rect 1871 8241 1927 8243
rect 2013 8241 2069 8243
rect 2155 8241 2211 8243
rect 2297 8241 2353 8243
rect 2439 8241 2495 8243
rect 25 8145 61 8155
rect 61 8145 81 8155
rect 167 8145 169 8155
rect 169 8145 221 8155
rect 221 8145 223 8155
rect 309 8145 329 8155
rect 329 8145 365 8155
rect 25 8099 81 8145
rect 167 8099 223 8145
rect 309 8099 365 8145
rect 451 8135 466 8155
rect 466 8135 507 8155
rect 593 8135 626 8155
rect 626 8135 649 8155
rect 735 8135 790 8155
rect 790 8135 791 8155
rect 877 8135 898 8155
rect 898 8135 933 8155
rect 1019 8135 1058 8155
rect 1058 8135 1075 8155
rect 1161 8135 1166 8155
rect 1166 8135 1217 8155
rect 1303 8135 1330 8155
rect 1330 8135 1359 8155
rect 1445 8135 1490 8155
rect 1490 8135 1501 8155
rect 1587 8135 1598 8155
rect 1598 8135 1643 8155
rect 1729 8135 1762 8155
rect 1762 8135 1785 8155
rect 1871 8135 1922 8155
rect 1922 8135 1927 8155
rect 2013 8135 2030 8155
rect 2030 8135 2069 8155
rect 2155 8135 2194 8155
rect 2194 8135 2211 8155
rect 2297 8135 2302 8155
rect 2302 8135 2353 8155
rect 2439 8135 2462 8155
rect 2462 8135 2495 8155
rect 451 8099 507 8135
rect 593 8099 649 8135
rect 735 8099 791 8135
rect 877 8099 933 8135
rect 1019 8099 1075 8135
rect 1161 8099 1217 8135
rect 1303 8099 1359 8135
rect 1445 8099 1501 8135
rect 1587 8099 1643 8135
rect 1729 8099 1785 8135
rect 1871 8099 1927 8135
rect 2013 8099 2069 8135
rect 2155 8099 2211 8135
rect 2297 8099 2353 8135
rect 2439 8099 2495 8135
rect 3403 8403 3459 8439
rect 3545 8403 3601 8439
rect 3687 8403 3743 8439
rect 3829 8403 3885 8439
rect 3971 8403 4027 8439
rect 4113 8403 4169 8439
rect 4255 8403 4311 8439
rect 4397 8403 4453 8439
rect 4539 8403 4595 8439
rect 4681 8403 4737 8439
rect 4823 8403 4879 8439
rect 4965 8403 5021 8439
rect 5107 8403 5163 8439
rect 5249 8403 5305 8439
rect 5391 8403 5447 8439
rect 3403 8383 3436 8403
rect 3436 8383 3459 8403
rect 3545 8383 3596 8403
rect 3596 8383 3601 8403
rect 3687 8383 3704 8403
rect 3704 8383 3743 8403
rect 3829 8383 3868 8403
rect 3868 8383 3885 8403
rect 3971 8383 3976 8403
rect 3976 8383 4027 8403
rect 4113 8383 4136 8403
rect 4136 8383 4169 8403
rect 4255 8383 4300 8403
rect 4300 8383 4311 8403
rect 4397 8383 4408 8403
rect 4408 8383 4453 8403
rect 4539 8383 4568 8403
rect 4568 8383 4595 8403
rect 4681 8383 4732 8403
rect 4732 8383 4737 8403
rect 4823 8383 4840 8403
rect 4840 8383 4879 8403
rect 4965 8383 5000 8403
rect 5000 8383 5021 8403
rect 5107 8383 5108 8403
rect 5108 8383 5163 8403
rect 5249 8383 5272 8403
rect 5272 8383 5305 8403
rect 5391 8383 5432 8403
rect 5432 8383 5447 8403
rect 5533 8413 5589 8439
rect 5675 8413 5731 8439
rect 5817 8413 5873 8439
rect 5533 8383 5569 8413
rect 5569 8383 5589 8413
rect 5675 8383 5677 8413
rect 5677 8383 5729 8413
rect 5729 8383 5731 8413
rect 5817 8383 5837 8413
rect 5837 8383 5873 8413
rect 3403 8295 3459 8297
rect 3545 8295 3601 8297
rect 3687 8295 3743 8297
rect 3829 8295 3885 8297
rect 3971 8295 4027 8297
rect 4113 8295 4169 8297
rect 4255 8295 4311 8297
rect 4397 8295 4453 8297
rect 4539 8295 4595 8297
rect 4681 8295 4737 8297
rect 4823 8295 4879 8297
rect 4965 8295 5021 8297
rect 5107 8295 5163 8297
rect 5249 8295 5305 8297
rect 5391 8295 5447 8297
rect 3403 8243 3436 8295
rect 3436 8243 3459 8295
rect 3545 8243 3596 8295
rect 3596 8243 3601 8295
rect 3687 8243 3704 8295
rect 3704 8243 3743 8295
rect 3829 8243 3868 8295
rect 3868 8243 3885 8295
rect 3971 8243 3976 8295
rect 3976 8243 4027 8295
rect 4113 8243 4136 8295
rect 4136 8243 4169 8295
rect 4255 8243 4300 8295
rect 4300 8243 4311 8295
rect 4397 8243 4408 8295
rect 4408 8243 4453 8295
rect 4539 8243 4568 8295
rect 4568 8243 4595 8295
rect 4681 8243 4732 8295
rect 4732 8243 4737 8295
rect 4823 8243 4840 8295
rect 4840 8243 4879 8295
rect 4965 8243 5000 8295
rect 5000 8243 5021 8295
rect 5107 8243 5108 8295
rect 5108 8243 5163 8295
rect 5249 8243 5272 8295
rect 5272 8243 5305 8295
rect 5391 8243 5432 8295
rect 5432 8243 5447 8295
rect 3403 8241 3459 8243
rect 3545 8241 3601 8243
rect 3687 8241 3743 8243
rect 3829 8241 3885 8243
rect 3971 8241 4027 8243
rect 4113 8241 4169 8243
rect 4255 8241 4311 8243
rect 4397 8241 4453 8243
rect 4539 8241 4595 8243
rect 4681 8241 4737 8243
rect 4823 8241 4879 8243
rect 4965 8241 5021 8243
rect 5107 8241 5163 8243
rect 5249 8241 5305 8243
rect 5391 8241 5447 8243
rect 5533 8253 5569 8297
rect 5569 8253 5589 8297
rect 5675 8253 5677 8297
rect 5677 8253 5729 8297
rect 5729 8253 5731 8297
rect 5817 8253 5837 8297
rect 5837 8253 5873 8297
rect 5533 8241 5589 8253
rect 5675 8241 5731 8253
rect 5817 8241 5873 8253
rect 3403 8135 3436 8155
rect 3436 8135 3459 8155
rect 3545 8135 3596 8155
rect 3596 8135 3601 8155
rect 3687 8135 3704 8155
rect 3704 8135 3743 8155
rect 3829 8135 3868 8155
rect 3868 8135 3885 8155
rect 3971 8135 3976 8155
rect 3976 8135 4027 8155
rect 4113 8135 4136 8155
rect 4136 8135 4169 8155
rect 4255 8135 4300 8155
rect 4300 8135 4311 8155
rect 4397 8135 4408 8155
rect 4408 8135 4453 8155
rect 4539 8135 4568 8155
rect 4568 8135 4595 8155
rect 4681 8135 4732 8155
rect 4732 8135 4737 8155
rect 4823 8135 4840 8155
rect 4840 8135 4879 8155
rect 4965 8135 5000 8155
rect 5000 8135 5021 8155
rect 5107 8135 5108 8155
rect 5108 8135 5163 8155
rect 5249 8135 5272 8155
rect 5272 8135 5305 8155
rect 5391 8135 5432 8155
rect 5432 8135 5447 8155
rect 3403 8099 3459 8135
rect 3545 8099 3601 8135
rect 3687 8099 3743 8135
rect 3829 8099 3885 8135
rect 3971 8099 4027 8135
rect 4113 8099 4169 8135
rect 4255 8099 4311 8135
rect 4397 8099 4453 8135
rect 4539 8099 4595 8135
rect 4681 8099 4737 8135
rect 4823 8099 4879 8135
rect 4965 8099 5021 8135
rect 5107 8099 5163 8135
rect 5249 8099 5305 8135
rect 5391 8099 5447 8135
rect 5533 8145 5569 8155
rect 5569 8145 5589 8155
rect 5675 8145 5677 8155
rect 5677 8145 5729 8155
rect 5729 8145 5731 8155
rect 5817 8145 5837 8155
rect 5837 8145 5873 8155
rect 5533 8099 5589 8145
rect 5675 8099 5731 8145
rect 5817 8099 5873 8145
rect 25 7821 61 7835
rect 61 7821 81 7835
rect 167 7821 169 7835
rect 169 7821 221 7835
rect 221 7821 223 7835
rect 309 7821 329 7835
rect 329 7821 365 7835
rect 25 7779 81 7821
rect 167 7779 223 7821
rect 309 7779 365 7821
rect 25 7657 81 7693
rect 167 7657 223 7693
rect 309 7657 365 7693
rect 25 7637 61 7657
rect 61 7637 81 7657
rect 167 7637 169 7657
rect 169 7637 221 7657
rect 221 7637 223 7657
rect 309 7637 329 7657
rect 329 7637 365 7657
rect 25 7549 81 7551
rect 167 7549 223 7551
rect 309 7549 365 7551
rect 25 7497 61 7549
rect 61 7497 81 7549
rect 167 7497 169 7549
rect 169 7497 221 7549
rect 221 7497 223 7549
rect 309 7497 329 7549
rect 329 7497 365 7549
rect 25 7495 81 7497
rect 167 7495 223 7497
rect 309 7495 365 7497
rect 25 7389 61 7409
rect 61 7389 81 7409
rect 167 7389 169 7409
rect 169 7389 221 7409
rect 221 7389 223 7409
rect 309 7389 329 7409
rect 329 7389 365 7409
rect 25 7353 81 7389
rect 167 7353 223 7389
rect 309 7353 365 7389
rect 25 7225 81 7267
rect 167 7225 223 7267
rect 309 7225 365 7267
rect 25 7211 61 7225
rect 61 7211 81 7225
rect 167 7211 169 7225
rect 169 7211 221 7225
rect 221 7211 223 7225
rect 309 7211 329 7225
rect 329 7211 365 7225
rect 5533 7821 5569 7835
rect 5569 7821 5589 7835
rect 5675 7821 5677 7835
rect 5677 7821 5729 7835
rect 5729 7821 5731 7835
rect 5817 7821 5837 7835
rect 5837 7821 5873 7835
rect 5533 7779 5589 7821
rect 5675 7779 5731 7821
rect 5817 7779 5873 7821
rect 5533 7657 5589 7693
rect 5675 7657 5731 7693
rect 5817 7657 5873 7693
rect 5533 7637 5569 7657
rect 5569 7637 5589 7657
rect 5675 7637 5677 7657
rect 5677 7637 5729 7657
rect 5729 7637 5731 7657
rect 5817 7637 5837 7657
rect 5837 7637 5873 7657
rect 5533 7549 5589 7551
rect 5675 7549 5731 7551
rect 5817 7549 5873 7551
rect 5533 7497 5569 7549
rect 5569 7497 5589 7549
rect 5675 7497 5677 7549
rect 5677 7497 5729 7549
rect 5729 7497 5731 7549
rect 5817 7497 5837 7549
rect 5837 7497 5873 7549
rect 5533 7495 5589 7497
rect 5675 7495 5731 7497
rect 5817 7495 5873 7497
rect 5533 7389 5569 7409
rect 5569 7389 5589 7409
rect 5675 7389 5677 7409
rect 5677 7389 5729 7409
rect 5729 7389 5731 7409
rect 5817 7389 5837 7409
rect 5837 7389 5873 7409
rect 5533 7353 5589 7389
rect 5675 7353 5731 7389
rect 5817 7353 5873 7389
rect 5533 7225 5589 7267
rect 5675 7225 5731 7267
rect 5817 7225 5873 7267
rect 5533 7211 5569 7225
rect 5569 7211 5589 7225
rect 5675 7211 5677 7225
rect 5677 7211 5729 7225
rect 5729 7211 5731 7225
rect 5817 7211 5837 7225
rect 5837 7211 5873 7225
rect 25 7117 81 7125
rect 167 7117 223 7125
rect 309 7117 365 7125
rect 25 7069 61 7117
rect 61 7069 81 7117
rect 167 7069 169 7117
rect 169 7069 221 7117
rect 221 7069 223 7117
rect 309 7069 329 7117
rect 329 7069 365 7117
rect 25 6957 61 6983
rect 61 6957 81 6983
rect 167 6957 169 6983
rect 169 6957 221 6983
rect 221 6957 223 6983
rect 309 6957 329 6983
rect 329 6957 365 6983
rect 25 6927 81 6957
rect 167 6927 223 6957
rect 309 6927 365 6957
rect 25 6793 81 6841
rect 167 6793 223 6841
rect 309 6793 365 6841
rect 25 6785 61 6793
rect 61 6785 81 6793
rect 167 6785 169 6793
rect 169 6785 221 6793
rect 221 6785 223 6793
rect 309 6785 329 6793
rect 329 6785 365 6793
rect 25 6685 81 6699
rect 167 6685 223 6699
rect 309 6685 365 6699
rect 25 6643 61 6685
rect 61 6643 81 6685
rect 167 6643 169 6685
rect 169 6643 221 6685
rect 221 6643 223 6685
rect 309 6643 329 6685
rect 329 6643 365 6685
rect 25 6525 61 6557
rect 61 6525 81 6557
rect 167 6525 169 6557
rect 169 6525 221 6557
rect 221 6525 223 6557
rect 309 6525 329 6557
rect 329 6525 365 6557
rect 25 6501 81 6525
rect 167 6501 223 6525
rect 309 6501 365 6525
rect 5533 7117 5589 7125
rect 5675 7117 5731 7125
rect 5817 7117 5873 7125
rect 5533 7069 5569 7117
rect 5569 7069 5589 7117
rect 5675 7069 5677 7117
rect 5677 7069 5729 7117
rect 5729 7069 5731 7117
rect 5817 7069 5837 7117
rect 5837 7069 5873 7117
rect 5533 6957 5569 6983
rect 5569 6957 5589 6983
rect 5675 6957 5677 6983
rect 5677 6957 5729 6983
rect 5729 6957 5731 6983
rect 5817 6957 5837 6983
rect 5837 6957 5873 6983
rect 5533 6927 5589 6957
rect 5675 6927 5731 6957
rect 5817 6927 5873 6957
rect 5533 6793 5589 6841
rect 5675 6793 5731 6841
rect 5817 6793 5873 6841
rect 5533 6785 5569 6793
rect 5569 6785 5589 6793
rect 5675 6785 5677 6793
rect 5677 6785 5729 6793
rect 5729 6785 5731 6793
rect 5817 6785 5837 6793
rect 5837 6785 5873 6793
rect 5533 6685 5589 6699
rect 5675 6685 5731 6699
rect 5817 6685 5873 6699
rect 5533 6643 5569 6685
rect 5569 6643 5589 6685
rect 5675 6643 5677 6685
rect 5677 6643 5729 6685
rect 5729 6643 5731 6685
rect 5817 6643 5837 6685
rect 5837 6643 5873 6685
rect 5533 6525 5569 6557
rect 5569 6525 5589 6557
rect 5675 6525 5677 6557
rect 5677 6525 5729 6557
rect 5729 6525 5731 6557
rect 5817 6525 5837 6557
rect 5837 6525 5873 6557
rect 5533 6501 5589 6525
rect 5675 6501 5731 6525
rect 5817 6501 5873 6525
rect 560 5656 579 5688
rect 579 5656 616 5688
rect 702 5656 739 5688
rect 739 5656 758 5688
rect 560 5632 616 5656
rect 702 5632 758 5656
rect 560 5492 616 5546
rect 702 5492 758 5546
rect 560 5490 579 5492
rect 579 5490 616 5492
rect 702 5490 739 5492
rect 739 5490 758 5492
rect 560 5384 616 5404
rect 702 5384 758 5404
rect 560 5348 579 5384
rect 579 5348 616 5384
rect 702 5348 739 5384
rect 739 5348 758 5384
rect 560 5224 579 5262
rect 579 5224 616 5262
rect 702 5224 739 5262
rect 739 5224 758 5262
rect 560 5206 616 5224
rect 702 5206 758 5224
rect 560 5116 579 5120
rect 579 5116 616 5120
rect 702 5116 739 5120
rect 739 5116 758 5120
rect 560 5064 616 5116
rect 702 5064 758 5116
rect 560 4952 616 4978
rect 702 4952 758 4978
rect 560 4922 579 4952
rect 579 4922 616 4952
rect 702 4922 739 4952
rect 739 4922 758 4952
rect 25 4611 81 4624
rect 167 4611 223 4624
rect 309 4611 365 4624
rect 25 4568 61 4611
rect 61 4568 81 4611
rect 167 4568 169 4611
rect 169 4568 221 4611
rect 221 4568 223 4611
rect 309 4568 329 4611
rect 329 4568 365 4611
rect 25 4451 61 4482
rect 61 4451 81 4482
rect 167 4451 169 4482
rect 169 4451 221 4482
rect 221 4451 223 4482
rect 309 4451 329 4482
rect 329 4451 365 4482
rect 25 4426 81 4451
rect 167 4426 223 4451
rect 309 4426 365 4451
rect 25 4287 81 4340
rect 167 4287 223 4340
rect 309 4287 365 4340
rect 25 4284 61 4287
rect 61 4284 81 4287
rect 167 4284 169 4287
rect 169 4284 221 4287
rect 221 4284 223 4287
rect 309 4284 329 4287
rect 329 4284 365 4287
rect 25 4179 81 4198
rect 167 4179 223 4198
rect 309 4179 365 4198
rect 25 4142 61 4179
rect 61 4142 81 4179
rect 167 4142 169 4179
rect 169 4142 221 4179
rect 221 4142 223 4179
rect 309 4142 329 4179
rect 329 4142 365 4179
rect 25 4019 61 4056
rect 61 4019 81 4056
rect 167 4019 169 4056
rect 169 4019 221 4056
rect 221 4019 223 4056
rect 309 4019 329 4056
rect 329 4019 365 4056
rect 25 4000 81 4019
rect 167 4000 223 4019
rect 309 4000 365 4019
rect 25 3911 61 3914
rect 61 3911 81 3914
rect 167 3911 169 3914
rect 169 3911 221 3914
rect 221 3911 223 3914
rect 309 3911 329 3914
rect 329 3911 365 3914
rect 25 3858 81 3911
rect 167 3858 223 3911
rect 309 3858 365 3911
rect 25 3747 81 3772
rect 167 3747 223 3772
rect 309 3747 365 3772
rect 25 3716 61 3747
rect 61 3716 81 3747
rect 167 3716 169 3747
rect 169 3716 221 3747
rect 221 3716 223 3747
rect 309 3716 329 3747
rect 329 3716 365 3747
rect 25 3587 61 3630
rect 61 3587 81 3630
rect 167 3587 169 3630
rect 169 3587 221 3630
rect 221 3587 223 3630
rect 309 3587 329 3630
rect 329 3587 365 3630
rect 25 3574 81 3587
rect 167 3574 223 3587
rect 309 3574 365 3587
rect 1508 5632 1564 5688
rect 1650 5632 1706 5688
rect 1792 5632 1848 5688
rect 1508 5490 1564 5546
rect 1650 5490 1706 5546
rect 1792 5490 1848 5546
rect 1508 5348 1564 5404
rect 1650 5348 1706 5404
rect 1792 5348 1848 5404
rect 1508 5206 1564 5262
rect 1650 5206 1706 5262
rect 1792 5206 1848 5262
rect 1508 5064 1564 5120
rect 1650 5064 1706 5120
rect 1792 5064 1848 5120
rect 1508 4922 1564 4978
rect 1650 4922 1706 4978
rect 1792 4922 1848 4978
rect 2520 5632 2576 5688
rect 2662 5632 2718 5688
rect 2804 5632 2860 5688
rect 2520 5490 2576 5546
rect 2662 5490 2718 5546
rect 2804 5490 2860 5546
rect 2520 5348 2576 5404
rect 2662 5348 2718 5404
rect 2804 5348 2860 5404
rect 2520 5206 2576 5262
rect 2662 5206 2718 5262
rect 2804 5206 2860 5262
rect 2520 5064 2576 5120
rect 2662 5064 2718 5120
rect 2804 5064 2860 5120
rect 2520 4922 2576 4978
rect 2662 4922 2718 4978
rect 2804 4922 2860 4978
rect 3038 5632 3094 5688
rect 3180 5632 3236 5688
rect 3322 5632 3378 5688
rect 3038 5490 3094 5546
rect 3180 5490 3236 5546
rect 3322 5490 3378 5546
rect 3038 5348 3094 5404
rect 3180 5348 3236 5404
rect 3322 5348 3378 5404
rect 3038 5206 3094 5262
rect 3180 5206 3236 5262
rect 3322 5206 3378 5262
rect 3038 5064 3094 5120
rect 3180 5064 3236 5120
rect 3322 5064 3378 5120
rect 3038 4922 3094 4978
rect 3180 4922 3236 4978
rect 3322 4922 3378 4978
rect 4050 5632 4106 5688
rect 4192 5632 4248 5688
rect 4334 5632 4390 5688
rect 4050 5490 4106 5546
rect 4192 5490 4248 5546
rect 4334 5490 4390 5546
rect 4050 5348 4106 5404
rect 4192 5348 4248 5404
rect 4334 5348 4390 5404
rect 4050 5206 4106 5262
rect 4192 5206 4248 5262
rect 4334 5206 4390 5262
rect 4050 5064 4106 5120
rect 4192 5064 4248 5120
rect 4334 5064 4390 5120
rect 4050 4922 4106 4978
rect 4192 4922 4248 4978
rect 4334 4922 4390 4978
rect 5140 5656 5159 5688
rect 5159 5656 5196 5688
rect 5282 5656 5319 5688
rect 5319 5656 5338 5688
rect 5140 5632 5196 5656
rect 5282 5632 5338 5656
rect 5140 5492 5196 5546
rect 5282 5492 5338 5546
rect 5140 5490 5159 5492
rect 5159 5490 5196 5492
rect 5282 5490 5319 5492
rect 5319 5490 5338 5492
rect 5140 5384 5196 5404
rect 5282 5384 5338 5404
rect 5140 5348 5159 5384
rect 5159 5348 5196 5384
rect 5282 5348 5319 5384
rect 5319 5348 5338 5384
rect 5140 5224 5159 5262
rect 5159 5224 5196 5262
rect 5282 5224 5319 5262
rect 5319 5224 5338 5262
rect 5140 5206 5196 5224
rect 5282 5206 5338 5224
rect 5140 5116 5159 5120
rect 5159 5116 5196 5120
rect 5282 5116 5319 5120
rect 5319 5116 5338 5120
rect 5140 5064 5196 5116
rect 5282 5064 5338 5116
rect 5140 4952 5196 4978
rect 5282 4952 5338 4978
rect 5140 4922 5159 4952
rect 5159 4922 5196 4952
rect 5282 4922 5319 4952
rect 5319 4922 5338 4952
rect 5533 4581 5569 4626
rect 5569 4581 5589 4626
rect 5675 4581 5677 4626
rect 5677 4581 5729 4626
rect 5729 4581 5731 4626
rect 5817 4581 5837 4626
rect 5837 4581 5873 4626
rect 5533 4570 5589 4581
rect 5675 4570 5731 4581
rect 5817 4570 5873 4581
rect 5533 4473 5569 4484
rect 5569 4473 5589 4484
rect 5675 4473 5677 4484
rect 5677 4473 5729 4484
rect 5729 4473 5731 4484
rect 5817 4473 5837 4484
rect 5837 4473 5873 4484
rect 5533 4428 5589 4473
rect 5675 4428 5731 4473
rect 5817 4428 5873 4473
rect 5533 4309 5589 4342
rect 5675 4309 5731 4342
rect 5817 4309 5873 4342
rect 5533 4286 5569 4309
rect 5569 4286 5589 4309
rect 5675 4286 5677 4309
rect 5677 4286 5729 4309
rect 5729 4286 5731 4309
rect 5817 4286 5837 4309
rect 5837 4286 5873 4309
rect 5533 4149 5569 4200
rect 5569 4149 5589 4200
rect 5675 4149 5677 4200
rect 5677 4149 5729 4200
rect 5729 4149 5731 4200
rect 5817 4149 5837 4200
rect 5837 4149 5873 4200
rect 5533 4144 5589 4149
rect 5675 4144 5731 4149
rect 5817 4144 5873 4149
rect 5533 4041 5569 4058
rect 5569 4041 5589 4058
rect 5675 4041 5677 4058
rect 5677 4041 5729 4058
rect 5729 4041 5731 4058
rect 5817 4041 5837 4058
rect 5837 4041 5873 4058
rect 5533 4002 5589 4041
rect 5675 4002 5731 4041
rect 5817 4002 5873 4041
rect 5533 3877 5589 3916
rect 5675 3877 5731 3916
rect 5817 3877 5873 3916
rect 5533 3860 5569 3877
rect 5569 3860 5589 3877
rect 5675 3860 5677 3877
rect 5677 3860 5729 3877
rect 5729 3860 5731 3877
rect 5817 3860 5837 3877
rect 5837 3860 5873 3877
rect 5533 3769 5589 3774
rect 5675 3769 5731 3774
rect 5817 3769 5873 3774
rect 5533 3718 5569 3769
rect 5569 3718 5589 3769
rect 5675 3718 5677 3769
rect 5677 3718 5729 3769
rect 5729 3718 5731 3769
rect 5817 3718 5837 3769
rect 5837 3718 5873 3769
rect 5533 3609 5569 3632
rect 5569 3609 5589 3632
rect 5675 3609 5677 3632
rect 5677 3609 5729 3632
rect 5729 3609 5731 3632
rect 5817 3609 5837 3632
rect 5837 3609 5873 3632
rect 5533 3576 5589 3609
rect 5675 3576 5731 3609
rect 5817 3576 5873 3609
rect 5533 3445 5589 3490
rect 5675 3445 5731 3490
rect 5817 3445 5873 3490
rect 5533 3434 5569 3445
rect 5569 3434 5589 3445
rect 5675 3434 5677 3445
rect 5677 3434 5729 3445
rect 5729 3434 5731 3445
rect 5817 3434 5837 3445
rect 5837 3434 5873 3445
rect 5533 3337 5589 3348
rect 5675 3337 5731 3348
rect 5817 3337 5873 3348
rect 5533 3292 5569 3337
rect 5569 3292 5589 3337
rect 5675 3292 5677 3337
rect 5677 3292 5729 3337
rect 5729 3292 5731 3337
rect 5817 3292 5837 3337
rect 5837 3292 5873 3337
rect 25 2769 61 2779
rect 61 2769 81 2779
rect 167 2769 169 2779
rect 169 2769 221 2779
rect 221 2769 223 2779
rect 309 2769 329 2779
rect 329 2769 365 2779
rect 25 2723 81 2769
rect 167 2723 223 2769
rect 309 2723 365 2769
rect 25 2605 81 2637
rect 167 2605 223 2637
rect 309 2605 365 2637
rect 25 2581 61 2605
rect 61 2581 81 2605
rect 167 2581 169 2605
rect 169 2581 221 2605
rect 221 2581 223 2605
rect 309 2581 329 2605
rect 329 2581 365 2605
rect 25 2445 61 2495
rect 61 2445 81 2495
rect 167 2445 169 2495
rect 169 2445 221 2495
rect 221 2445 223 2495
rect 309 2445 329 2495
rect 329 2445 365 2495
rect 25 2439 81 2445
rect 167 2439 223 2445
rect 309 2439 365 2445
rect 25 2337 61 2353
rect 61 2337 81 2353
rect 167 2337 169 2353
rect 169 2337 221 2353
rect 221 2337 223 2353
rect 309 2337 329 2353
rect 329 2337 365 2353
rect 25 2297 81 2337
rect 167 2297 223 2337
rect 309 2297 365 2337
rect 25 2173 81 2211
rect 167 2173 223 2211
rect 309 2173 365 2211
rect 25 2155 61 2173
rect 61 2155 81 2173
rect 167 2155 169 2173
rect 169 2155 221 2173
rect 221 2155 223 2173
rect 309 2155 329 2173
rect 329 2155 365 2173
rect 25 2065 81 2069
rect 167 2065 223 2069
rect 309 2065 365 2069
rect 25 2013 61 2065
rect 61 2013 81 2065
rect 167 2013 169 2065
rect 169 2013 221 2065
rect 221 2013 223 2065
rect 309 2013 329 2065
rect 329 2013 365 2065
rect 25 1905 61 1927
rect 61 1905 81 1927
rect 167 1905 169 1927
rect 169 1905 221 1927
rect 221 1905 223 1927
rect 309 1905 329 1927
rect 329 1905 365 1927
rect 25 1871 81 1905
rect 167 1871 223 1905
rect 309 1871 365 1905
rect 25 1741 81 1785
rect 167 1741 223 1785
rect 309 1741 365 1785
rect 25 1729 61 1741
rect 61 1729 81 1741
rect 167 1729 169 1741
rect 169 1729 221 1741
rect 221 1729 223 1741
rect 309 1729 329 1741
rect 329 1729 365 1741
rect 560 1416 616 1418
rect 702 1416 758 1418
rect 560 1364 579 1416
rect 579 1364 616 1416
rect 702 1364 739 1416
rect 739 1364 758 1416
rect 560 1362 616 1364
rect 702 1362 758 1364
rect 560 1256 579 1276
rect 579 1256 616 1276
rect 702 1256 739 1276
rect 739 1256 758 1276
rect 560 1220 616 1256
rect 702 1220 758 1256
rect 560 1092 616 1134
rect 702 1092 758 1134
rect 560 1078 579 1092
rect 579 1078 616 1092
rect 702 1078 739 1092
rect 739 1078 758 1092
rect 560 984 616 992
rect 702 984 758 992
rect 560 936 579 984
rect 579 936 616 984
rect 702 936 739 984
rect 739 936 758 984
rect 1508 1415 1564 1418
rect 1650 1415 1706 1418
rect 1792 1415 1848 1418
rect 1508 1362 1564 1415
rect 1650 1362 1706 1415
rect 1792 1362 1848 1415
rect 1508 1220 1564 1276
rect 1650 1220 1706 1276
rect 1792 1220 1848 1276
rect 1508 1078 1564 1134
rect 1650 1078 1706 1134
rect 1792 1078 1848 1134
rect 1508 936 1564 992
rect 1650 936 1706 992
rect 1792 936 1848 992
rect 2535 1415 2554 1418
rect 2554 1415 2591 1418
rect 2677 1415 2710 1418
rect 2710 1415 2733 1418
rect 2535 1362 2591 1415
rect 2677 1362 2733 1415
rect 2535 1220 2591 1276
rect 2677 1220 2733 1276
rect 2535 1078 2591 1134
rect 2677 1078 2733 1134
rect 2535 936 2591 992
rect 2677 936 2733 992
rect 3166 1415 3185 1418
rect 3185 1415 3222 1418
rect 3308 1415 3341 1418
rect 3341 1415 3364 1418
rect 3166 1362 3222 1415
rect 3308 1362 3364 1415
rect 3166 1220 3222 1276
rect 3308 1220 3364 1276
rect 3166 1078 3222 1134
rect 3308 1078 3364 1134
rect 3166 936 3222 992
rect 3308 936 3364 992
rect 4050 1415 4106 1418
rect 4192 1415 4248 1418
rect 4334 1415 4390 1418
rect 4050 1362 4106 1415
rect 4192 1362 4248 1415
rect 4334 1362 4390 1415
rect 4050 1220 4106 1276
rect 4192 1220 4248 1276
rect 4334 1220 4390 1276
rect 4050 1078 4106 1134
rect 4192 1078 4248 1134
rect 4334 1078 4390 1134
rect 4050 936 4106 992
rect 4192 936 4248 992
rect 4334 936 4390 992
rect 5533 2981 5569 3033
rect 5569 2981 5589 3033
rect 5675 2981 5677 3033
rect 5677 2981 5729 3033
rect 5729 2981 5731 3033
rect 5817 2981 5837 3033
rect 5837 2981 5873 3033
rect 5533 2977 5589 2981
rect 5675 2977 5731 2981
rect 5817 2977 5873 2981
rect 5533 2873 5569 2891
rect 5569 2873 5589 2891
rect 5675 2873 5677 2891
rect 5677 2873 5729 2891
rect 5729 2873 5731 2891
rect 5817 2873 5837 2891
rect 5837 2873 5873 2891
rect 5533 2835 5589 2873
rect 5675 2835 5731 2873
rect 5817 2835 5873 2873
rect 5533 2709 5589 2749
rect 5675 2709 5731 2749
rect 5817 2709 5873 2749
rect 5533 2693 5569 2709
rect 5569 2693 5589 2709
rect 5675 2693 5677 2709
rect 5677 2693 5729 2709
rect 5729 2693 5731 2709
rect 5817 2693 5837 2709
rect 5837 2693 5873 2709
rect 5533 2601 5589 2607
rect 5675 2601 5731 2607
rect 5817 2601 5873 2607
rect 5533 2551 5569 2601
rect 5569 2551 5589 2601
rect 5675 2551 5677 2601
rect 5677 2551 5729 2601
rect 5729 2551 5731 2601
rect 5817 2551 5837 2601
rect 5837 2551 5873 2601
rect 5533 2441 5569 2465
rect 5569 2441 5589 2465
rect 5675 2441 5677 2465
rect 5677 2441 5729 2465
rect 5729 2441 5731 2465
rect 5817 2441 5837 2465
rect 5837 2441 5873 2465
rect 5533 2409 5589 2441
rect 5675 2409 5731 2441
rect 5817 2409 5873 2441
rect 5533 2277 5589 2323
rect 5675 2277 5731 2323
rect 5817 2277 5873 2323
rect 5533 2267 5569 2277
rect 5569 2267 5589 2277
rect 5675 2267 5677 2277
rect 5677 2267 5729 2277
rect 5729 2267 5731 2277
rect 5817 2267 5837 2277
rect 5837 2267 5873 2277
rect 5533 2169 5589 2181
rect 5675 2169 5731 2181
rect 5817 2169 5873 2181
rect 5533 2125 5569 2169
rect 5569 2125 5589 2169
rect 5675 2125 5677 2169
rect 5677 2125 5729 2169
rect 5729 2125 5731 2169
rect 5817 2125 5837 2169
rect 5837 2125 5873 2169
rect 5533 2009 5569 2039
rect 5569 2009 5589 2039
rect 5675 2009 5677 2039
rect 5677 2009 5729 2039
rect 5729 2009 5731 2039
rect 5817 2009 5837 2039
rect 5837 2009 5873 2039
rect 5533 1983 5589 2009
rect 5675 1983 5731 2009
rect 5817 1983 5873 2009
rect 5533 1845 5589 1897
rect 5675 1845 5731 1897
rect 5817 1845 5873 1897
rect 5533 1841 5569 1845
rect 5569 1841 5589 1845
rect 5675 1841 5677 1845
rect 5677 1841 5729 1845
rect 5729 1841 5731 1845
rect 5817 1841 5837 1845
rect 5837 1841 5873 1845
rect 5533 1737 5589 1755
rect 5675 1737 5731 1755
rect 5817 1737 5873 1755
rect 5533 1699 5569 1737
rect 5569 1699 5589 1737
rect 5675 1699 5677 1737
rect 5677 1699 5729 1737
rect 5729 1699 5731 1737
rect 5817 1699 5837 1737
rect 5837 1699 5873 1737
rect 5140 1416 5196 1418
rect 5282 1416 5338 1418
rect 5140 1364 5159 1416
rect 5159 1364 5196 1416
rect 5282 1364 5319 1416
rect 5319 1364 5338 1416
rect 5140 1362 5196 1364
rect 5282 1362 5338 1364
rect 5140 1256 5159 1276
rect 5159 1256 5196 1276
rect 5282 1256 5319 1276
rect 5319 1256 5338 1276
rect 5140 1220 5196 1256
rect 5282 1220 5338 1256
rect 5140 1092 5196 1134
rect 5282 1092 5338 1134
rect 5140 1078 5159 1092
rect 5159 1078 5196 1092
rect 5282 1078 5319 1092
rect 5319 1078 5338 1092
rect 5140 984 5196 992
rect 5282 984 5338 992
rect 5140 936 5159 984
rect 5159 936 5196 984
rect 5282 936 5319 984
rect 5319 936 5338 984
rect 578 768 634 787
rect 720 768 776 787
rect 862 768 918 787
rect 1004 768 1060 787
rect 1146 768 1202 787
rect 1288 768 1344 787
rect 1430 768 1486 787
rect 1572 768 1628 787
rect 1714 768 1770 787
rect 1856 768 1912 787
rect 1998 768 2054 787
rect 2140 768 2196 787
rect 2282 768 2338 787
rect 2424 768 2480 787
rect 2566 768 2622 787
rect 578 731 579 768
rect 579 731 631 768
rect 631 731 634 768
rect 720 731 739 768
rect 739 731 776 768
rect 862 731 869 768
rect 869 731 918 768
rect 1004 731 1033 768
rect 1033 731 1060 768
rect 1146 731 1193 768
rect 1193 731 1202 768
rect 1288 731 1301 768
rect 1301 731 1344 768
rect 1430 731 1465 768
rect 1465 731 1486 768
rect 1572 731 1573 768
rect 1573 731 1625 768
rect 1625 731 1628 768
rect 1714 731 1733 768
rect 1733 731 1770 768
rect 1856 731 1897 768
rect 1897 731 1912 768
rect 1998 731 2005 768
rect 2005 731 2054 768
rect 2140 731 2165 768
rect 2165 731 2196 768
rect 2282 731 2329 768
rect 2329 731 2338 768
rect 2424 731 2437 768
rect 2437 731 2480 768
rect 2566 731 2597 768
rect 2597 731 2622 768
rect 2708 731 2764 787
rect 578 608 579 645
rect 579 608 631 645
rect 631 608 634 645
rect 720 608 739 645
rect 739 608 776 645
rect 862 608 869 645
rect 869 608 918 645
rect 1004 608 1033 645
rect 1033 608 1060 645
rect 1146 608 1193 645
rect 1193 608 1202 645
rect 1288 608 1301 645
rect 1301 608 1344 645
rect 1430 608 1465 645
rect 1465 608 1486 645
rect 1572 608 1573 645
rect 1573 608 1625 645
rect 1625 608 1628 645
rect 1714 608 1733 645
rect 1733 608 1770 645
rect 1856 608 1897 645
rect 1897 608 1912 645
rect 1998 608 2005 645
rect 2005 608 2054 645
rect 2140 608 2165 645
rect 2165 608 2196 645
rect 2282 608 2329 645
rect 2329 608 2338 645
rect 2424 608 2437 645
rect 2437 608 2480 645
rect 2566 608 2597 645
rect 2597 608 2622 645
rect 578 589 634 608
rect 720 589 776 608
rect 862 589 918 608
rect 1004 589 1060 608
rect 1146 589 1202 608
rect 1288 589 1344 608
rect 1430 589 1486 608
rect 1572 589 1628 608
rect 1714 589 1770 608
rect 1856 589 1912 608
rect 1998 589 2054 608
rect 2140 589 2196 608
rect 2282 589 2338 608
rect 2424 589 2480 608
rect 2566 589 2622 608
rect 2708 589 2764 645
rect 3134 731 3190 787
rect 3276 768 3332 787
rect 3418 768 3474 787
rect 3560 768 3616 787
rect 3702 768 3758 787
rect 3844 768 3900 787
rect 3986 768 4042 787
rect 4128 768 4184 787
rect 4270 768 4326 787
rect 4412 768 4468 787
rect 4554 768 4610 787
rect 4696 768 4752 787
rect 4838 768 4894 787
rect 4980 768 5036 787
rect 5122 768 5178 787
rect 5264 768 5320 787
rect 3276 731 3301 768
rect 3301 731 3332 768
rect 3418 731 3461 768
rect 3461 731 3474 768
rect 3560 731 3569 768
rect 3569 731 3616 768
rect 3702 731 3733 768
rect 3733 731 3758 768
rect 3844 731 3893 768
rect 3893 731 3900 768
rect 3986 731 4001 768
rect 4001 731 4042 768
rect 4128 731 4165 768
rect 4165 731 4184 768
rect 4270 731 4273 768
rect 4273 731 4325 768
rect 4325 731 4326 768
rect 4412 731 4433 768
rect 4433 731 4468 768
rect 4554 731 4597 768
rect 4597 731 4610 768
rect 4696 731 4705 768
rect 4705 731 4752 768
rect 4838 731 4865 768
rect 4865 731 4894 768
rect 4980 731 5029 768
rect 5029 731 5036 768
rect 5122 731 5159 768
rect 5159 731 5178 768
rect 5264 731 5267 768
rect 5267 731 5319 768
rect 5319 731 5320 768
rect 3134 589 3190 645
rect 3276 608 3301 645
rect 3301 608 3332 645
rect 3418 608 3461 645
rect 3461 608 3474 645
rect 3560 608 3569 645
rect 3569 608 3616 645
rect 3702 608 3733 645
rect 3733 608 3758 645
rect 3844 608 3893 645
rect 3893 608 3900 645
rect 3986 608 4001 645
rect 4001 608 4042 645
rect 4128 608 4165 645
rect 4165 608 4184 645
rect 4270 608 4273 645
rect 4273 608 4325 645
rect 4325 608 4326 645
rect 4412 608 4433 645
rect 4433 608 4468 645
rect 4554 608 4597 645
rect 4597 608 4610 645
rect 4696 608 4705 645
rect 4705 608 4752 645
rect 4838 608 4865 645
rect 4865 608 4894 645
rect 4980 608 5029 645
rect 5029 608 5036 645
rect 5122 608 5159 645
rect 5159 608 5178 645
rect 5264 608 5267 645
rect 5267 608 5319 645
rect 5319 608 5320 645
rect 3276 589 3332 608
rect 3418 589 3474 608
rect 3560 589 3616 608
rect 3702 589 3758 608
rect 3844 589 3900 608
rect 3986 589 4042 608
rect 4128 589 4184 608
rect 4270 589 4326 608
rect 4412 589 4468 608
rect 4554 589 4610 608
rect 4696 589 4752 608
rect 4838 589 4894 608
rect 4980 589 5036 608
rect 5122 589 5178 608
rect 5264 589 5320 608
<< metal3 >>
rect 15 8439 2505 8449
rect 15 8383 25 8439
rect 81 8383 167 8439
rect 223 8383 309 8439
rect 365 8383 451 8439
rect 507 8383 593 8439
rect 649 8383 735 8439
rect 791 8383 877 8439
rect 933 8383 1019 8439
rect 1075 8383 1161 8439
rect 1217 8383 1303 8439
rect 1359 8383 1445 8439
rect 1501 8383 1587 8439
rect 1643 8383 1729 8439
rect 1785 8383 1871 8439
rect 1927 8383 2013 8439
rect 2069 8383 2155 8439
rect 2211 8383 2297 8439
rect 2353 8383 2439 8439
rect 2495 8383 2505 8439
rect 15 8297 2505 8383
rect 15 8241 25 8297
rect 81 8241 167 8297
rect 223 8241 309 8297
rect 365 8241 451 8297
rect 507 8241 593 8297
rect 649 8241 735 8297
rect 791 8241 877 8297
rect 933 8241 1019 8297
rect 1075 8241 1161 8297
rect 1217 8241 1303 8297
rect 1359 8241 1445 8297
rect 1501 8241 1587 8297
rect 1643 8241 1729 8297
rect 1785 8241 1871 8297
rect 1927 8241 2013 8297
rect 2069 8241 2155 8297
rect 2211 8241 2297 8297
rect 2353 8241 2439 8297
rect 2495 8241 2505 8297
rect 15 8155 2505 8241
rect 15 8099 25 8155
rect 81 8099 167 8155
rect 223 8099 309 8155
rect 365 8099 451 8155
rect 507 8099 593 8155
rect 649 8099 735 8155
rect 791 8099 877 8155
rect 933 8099 1019 8155
rect 1075 8099 1161 8155
rect 1217 8099 1303 8155
rect 1359 8099 1445 8155
rect 1501 8099 1587 8155
rect 1643 8099 1729 8155
rect 1785 8099 1871 8155
rect 1927 8099 2013 8155
rect 2069 8099 2155 8155
rect 2211 8099 2297 8155
rect 2353 8099 2439 8155
rect 2495 8099 2505 8155
rect 15 8089 2505 8099
rect 3393 8439 5883 8449
rect 3393 8383 3403 8439
rect 3459 8383 3545 8439
rect 3601 8383 3687 8439
rect 3743 8383 3829 8439
rect 3885 8383 3971 8439
rect 4027 8383 4113 8439
rect 4169 8383 4255 8439
rect 4311 8383 4397 8439
rect 4453 8383 4539 8439
rect 4595 8383 4681 8439
rect 4737 8383 4823 8439
rect 4879 8383 4965 8439
rect 5021 8383 5107 8439
rect 5163 8383 5249 8439
rect 5305 8383 5391 8439
rect 5447 8383 5533 8439
rect 5589 8383 5675 8439
rect 5731 8383 5817 8439
rect 5873 8383 5883 8439
rect 3393 8297 5883 8383
rect 3393 8241 3403 8297
rect 3459 8241 3545 8297
rect 3601 8241 3687 8297
rect 3743 8241 3829 8297
rect 3885 8241 3971 8297
rect 4027 8241 4113 8297
rect 4169 8241 4255 8297
rect 4311 8241 4397 8297
rect 4453 8241 4539 8297
rect 4595 8241 4681 8297
rect 4737 8241 4823 8297
rect 4879 8241 4965 8297
rect 5021 8241 5107 8297
rect 5163 8241 5249 8297
rect 5305 8241 5391 8297
rect 5447 8241 5533 8297
rect 5589 8241 5675 8297
rect 5731 8241 5817 8297
rect 5873 8241 5883 8297
rect 3393 8155 5883 8241
rect 3393 8099 3403 8155
rect 3459 8099 3545 8155
rect 3601 8099 3687 8155
rect 3743 8099 3829 8155
rect 3885 8099 3971 8155
rect 4027 8099 4113 8155
rect 4169 8099 4255 8155
rect 4311 8099 4397 8155
rect 4453 8099 4539 8155
rect 4595 8099 4681 8155
rect 4737 8099 4823 8155
rect 4879 8099 4965 8155
rect 5021 8099 5107 8155
rect 5163 8099 5249 8155
rect 5305 8099 5391 8155
rect 5447 8099 5533 8155
rect 5589 8099 5675 8155
rect 5731 8099 5817 8155
rect 5873 8099 5883 8155
rect 3393 8089 5883 8099
rect 15 7835 375 7845
rect 15 7779 25 7835
rect 81 7779 167 7835
rect 223 7779 309 7835
rect 365 7779 375 7835
rect 15 7693 375 7779
rect 15 7637 25 7693
rect 81 7637 167 7693
rect 223 7637 309 7693
rect 365 7637 375 7693
rect 15 7551 375 7637
rect 15 7495 25 7551
rect 81 7495 167 7551
rect 223 7495 309 7551
rect 365 7495 375 7551
rect 15 7409 375 7495
rect 15 7353 25 7409
rect 81 7353 167 7409
rect 223 7353 309 7409
rect 365 7353 375 7409
rect 15 7267 375 7353
rect 15 7211 25 7267
rect 81 7211 167 7267
rect 223 7211 309 7267
rect 365 7211 375 7267
rect 15 7125 375 7211
rect 15 7069 25 7125
rect 81 7069 167 7125
rect 223 7069 309 7125
rect 365 7069 375 7125
rect 15 6983 375 7069
rect 15 6927 25 6983
rect 81 6927 167 6983
rect 223 6927 309 6983
rect 365 6927 375 6983
rect 15 6841 375 6927
rect 15 6785 25 6841
rect 81 6785 167 6841
rect 223 6785 309 6841
rect 365 6785 375 6841
rect 15 6699 375 6785
rect 15 6643 25 6699
rect 81 6643 167 6699
rect 223 6643 309 6699
rect 365 6643 375 6699
rect 15 6557 375 6643
rect 15 6501 25 6557
rect 81 6501 167 6557
rect 223 6501 309 6557
rect 365 6501 375 6557
rect 15 6491 375 6501
rect 5523 7835 5883 7845
rect 5523 7779 5533 7835
rect 5589 7779 5675 7835
rect 5731 7779 5817 7835
rect 5873 7779 5883 7835
rect 5523 7693 5883 7779
rect 5523 7637 5533 7693
rect 5589 7637 5675 7693
rect 5731 7637 5817 7693
rect 5873 7637 5883 7693
rect 5523 7551 5883 7637
rect 5523 7495 5533 7551
rect 5589 7495 5675 7551
rect 5731 7495 5817 7551
rect 5873 7495 5883 7551
rect 5523 7409 5883 7495
rect 5523 7353 5533 7409
rect 5589 7353 5675 7409
rect 5731 7353 5817 7409
rect 5873 7353 5883 7409
rect 5523 7267 5883 7353
rect 5523 7211 5533 7267
rect 5589 7211 5675 7267
rect 5731 7211 5817 7267
rect 5873 7211 5883 7267
rect 5523 7125 5883 7211
rect 5523 7069 5533 7125
rect 5589 7069 5675 7125
rect 5731 7069 5817 7125
rect 5873 7069 5883 7125
rect 5523 6983 5883 7069
rect 5523 6927 5533 6983
rect 5589 6927 5675 6983
rect 5731 6927 5817 6983
rect 5873 6927 5883 6983
rect 5523 6841 5883 6927
rect 5523 6785 5533 6841
rect 5589 6785 5675 6841
rect 5731 6785 5817 6841
rect 5873 6785 5883 6841
rect 5523 6699 5883 6785
rect 5523 6643 5533 6699
rect 5589 6643 5675 6699
rect 5731 6643 5817 6699
rect 5873 6643 5883 6699
rect 5523 6557 5883 6643
rect 5523 6501 5533 6557
rect 5589 6501 5675 6557
rect 5731 6501 5817 6557
rect 5873 6501 5883 6557
rect 5523 6491 5883 6501
rect 550 5688 768 5698
rect 550 5632 560 5688
rect 616 5632 702 5688
rect 758 5632 768 5688
rect 550 5546 768 5632
rect 550 5490 560 5546
rect 616 5490 702 5546
rect 758 5490 768 5546
rect 550 5404 768 5490
rect 550 5348 560 5404
rect 616 5348 702 5404
rect 758 5348 768 5404
rect 550 5262 768 5348
rect 550 5206 560 5262
rect 616 5206 702 5262
rect 758 5206 768 5262
rect 550 5120 768 5206
rect 550 5064 560 5120
rect 616 5064 702 5120
rect 758 5064 768 5120
rect 550 4978 768 5064
rect 550 4922 560 4978
rect 616 4922 702 4978
rect 758 4922 768 4978
rect 550 4912 768 4922
rect 1498 5688 1858 5698
rect 1498 5632 1508 5688
rect 1564 5632 1650 5688
rect 1706 5632 1792 5688
rect 1848 5632 1858 5688
rect 1498 5546 1858 5632
rect 1498 5490 1508 5546
rect 1564 5490 1650 5546
rect 1706 5490 1792 5546
rect 1848 5490 1858 5546
rect 1498 5404 1858 5490
rect 1498 5348 1508 5404
rect 1564 5348 1650 5404
rect 1706 5348 1792 5404
rect 1848 5348 1858 5404
rect 1498 5262 1858 5348
rect 1498 5206 1508 5262
rect 1564 5206 1650 5262
rect 1706 5206 1792 5262
rect 1848 5206 1858 5262
rect 1498 5120 1858 5206
rect 1498 5064 1508 5120
rect 1564 5064 1650 5120
rect 1706 5064 1792 5120
rect 1848 5064 1858 5120
rect 1498 4978 1858 5064
rect 1498 4922 1508 4978
rect 1564 4922 1650 4978
rect 1706 4922 1792 4978
rect 1848 4922 1858 4978
rect 1498 4912 1858 4922
rect 2510 5688 2870 5698
rect 2510 5632 2520 5688
rect 2576 5632 2662 5688
rect 2718 5632 2804 5688
rect 2860 5632 2870 5688
rect 2510 5546 2870 5632
rect 2510 5490 2520 5546
rect 2576 5490 2662 5546
rect 2718 5490 2804 5546
rect 2860 5490 2870 5546
rect 2510 5404 2870 5490
rect 2510 5348 2520 5404
rect 2576 5348 2662 5404
rect 2718 5348 2804 5404
rect 2860 5348 2870 5404
rect 2510 5262 2870 5348
rect 2510 5206 2520 5262
rect 2576 5206 2662 5262
rect 2718 5206 2804 5262
rect 2860 5206 2870 5262
rect 2510 5120 2870 5206
rect 2510 5064 2520 5120
rect 2576 5064 2662 5120
rect 2718 5064 2804 5120
rect 2860 5064 2870 5120
rect 2510 4978 2870 5064
rect 2510 4922 2520 4978
rect 2576 4922 2662 4978
rect 2718 4922 2804 4978
rect 2860 4922 2870 4978
rect 2510 4912 2870 4922
rect 3028 5688 3388 5698
rect 3028 5632 3038 5688
rect 3094 5632 3180 5688
rect 3236 5632 3322 5688
rect 3378 5632 3388 5688
rect 3028 5546 3388 5632
rect 3028 5490 3038 5546
rect 3094 5490 3180 5546
rect 3236 5490 3322 5546
rect 3378 5490 3388 5546
rect 3028 5404 3388 5490
rect 3028 5348 3038 5404
rect 3094 5348 3180 5404
rect 3236 5348 3322 5404
rect 3378 5348 3388 5404
rect 3028 5262 3388 5348
rect 3028 5206 3038 5262
rect 3094 5206 3180 5262
rect 3236 5206 3322 5262
rect 3378 5206 3388 5262
rect 3028 5120 3388 5206
rect 3028 5064 3038 5120
rect 3094 5064 3180 5120
rect 3236 5064 3322 5120
rect 3378 5064 3388 5120
rect 3028 4978 3388 5064
rect 3028 4922 3038 4978
rect 3094 4922 3180 4978
rect 3236 4922 3322 4978
rect 3378 4922 3388 4978
rect 3028 4912 3388 4922
rect 4040 5688 4400 5698
rect 4040 5632 4050 5688
rect 4106 5632 4192 5688
rect 4248 5632 4334 5688
rect 4390 5632 4400 5688
rect 4040 5546 4400 5632
rect 4040 5490 4050 5546
rect 4106 5490 4192 5546
rect 4248 5490 4334 5546
rect 4390 5490 4400 5546
rect 4040 5404 4400 5490
rect 4040 5348 4050 5404
rect 4106 5348 4192 5404
rect 4248 5348 4334 5404
rect 4390 5348 4400 5404
rect 4040 5262 4400 5348
rect 4040 5206 4050 5262
rect 4106 5206 4192 5262
rect 4248 5206 4334 5262
rect 4390 5206 4400 5262
rect 4040 5120 4400 5206
rect 4040 5064 4050 5120
rect 4106 5064 4192 5120
rect 4248 5064 4334 5120
rect 4390 5064 4400 5120
rect 4040 4978 4400 5064
rect 4040 4922 4050 4978
rect 4106 4922 4192 4978
rect 4248 4922 4334 4978
rect 4390 4922 4400 4978
rect 4040 4912 4400 4922
rect 5130 5688 5348 5698
rect 5130 5632 5140 5688
rect 5196 5632 5282 5688
rect 5338 5632 5348 5688
rect 5130 5546 5348 5632
rect 5130 5490 5140 5546
rect 5196 5490 5282 5546
rect 5338 5490 5348 5546
rect 5130 5404 5348 5490
rect 5130 5348 5140 5404
rect 5196 5348 5282 5404
rect 5338 5348 5348 5404
rect 5130 5262 5348 5348
rect 5130 5206 5140 5262
rect 5196 5206 5282 5262
rect 5338 5206 5348 5262
rect 5130 5120 5348 5206
rect 5130 5064 5140 5120
rect 5196 5064 5282 5120
rect 5338 5064 5348 5120
rect 5130 4978 5348 5064
rect 5130 4922 5140 4978
rect 5196 4922 5282 4978
rect 5338 4922 5348 4978
rect 5130 4912 5348 4922
rect 15 4624 375 4634
rect 15 4568 25 4624
rect 81 4568 167 4624
rect 223 4568 309 4624
rect 365 4568 375 4624
rect 15 4482 375 4568
rect 15 4426 25 4482
rect 81 4426 167 4482
rect 223 4426 309 4482
rect 365 4426 375 4482
rect 15 4340 375 4426
rect 15 4284 25 4340
rect 81 4284 167 4340
rect 223 4284 309 4340
rect 365 4284 375 4340
rect 15 4198 375 4284
rect 15 4142 25 4198
rect 81 4142 167 4198
rect 223 4142 309 4198
rect 365 4142 375 4198
rect 15 4056 375 4142
rect 15 4000 25 4056
rect 81 4000 167 4056
rect 223 4000 309 4056
rect 365 4000 375 4056
rect 15 3914 375 4000
rect 15 3858 25 3914
rect 81 3858 167 3914
rect 223 3858 309 3914
rect 365 3858 375 3914
rect 15 3772 375 3858
rect 15 3716 25 3772
rect 81 3716 167 3772
rect 223 3716 309 3772
rect 365 3716 375 3772
rect 15 3630 375 3716
rect 15 3574 25 3630
rect 81 3574 167 3630
rect 223 3574 309 3630
rect 365 3574 375 3630
rect 15 3564 375 3574
rect 5523 4626 5883 4636
rect 5523 4570 5533 4626
rect 5589 4570 5675 4626
rect 5731 4570 5817 4626
rect 5873 4570 5883 4626
rect 5523 4484 5883 4570
rect 5523 4428 5533 4484
rect 5589 4428 5675 4484
rect 5731 4428 5817 4484
rect 5873 4428 5883 4484
rect 5523 4342 5883 4428
rect 5523 4286 5533 4342
rect 5589 4286 5675 4342
rect 5731 4286 5817 4342
rect 5873 4286 5883 4342
rect 5523 4200 5883 4286
rect 5523 4144 5533 4200
rect 5589 4144 5675 4200
rect 5731 4144 5817 4200
rect 5873 4144 5883 4200
rect 5523 4058 5883 4144
rect 5523 4002 5533 4058
rect 5589 4002 5675 4058
rect 5731 4002 5817 4058
rect 5873 4002 5883 4058
rect 5523 3916 5883 4002
rect 5523 3860 5533 3916
rect 5589 3860 5675 3916
rect 5731 3860 5817 3916
rect 5873 3860 5883 3916
rect 5523 3774 5883 3860
rect 5523 3718 5533 3774
rect 5589 3718 5675 3774
rect 5731 3718 5817 3774
rect 5873 3718 5883 3774
rect 5523 3632 5883 3718
rect 5523 3576 5533 3632
rect 5589 3576 5675 3632
rect 5731 3576 5817 3632
rect 5873 3576 5883 3632
rect 5523 3490 5883 3576
rect 5523 3434 5533 3490
rect 5589 3434 5675 3490
rect 5731 3434 5817 3490
rect 5873 3434 5883 3490
rect 5523 3348 5883 3434
rect 5523 3292 5533 3348
rect 5589 3292 5675 3348
rect 5731 3292 5817 3348
rect 5873 3292 5883 3348
rect 5523 3282 5883 3292
rect 5523 3033 5883 3043
rect 5523 2977 5533 3033
rect 5589 2977 5675 3033
rect 5731 2977 5817 3033
rect 5873 2977 5883 3033
rect 5523 2891 5883 2977
rect 5523 2835 5533 2891
rect 5589 2835 5675 2891
rect 5731 2835 5817 2891
rect 5873 2835 5883 2891
rect 15 2779 375 2789
rect 15 2723 25 2779
rect 81 2723 167 2779
rect 223 2723 309 2779
rect 365 2723 375 2779
rect 15 2637 375 2723
rect 15 2581 25 2637
rect 81 2581 167 2637
rect 223 2581 309 2637
rect 365 2581 375 2637
rect 15 2495 375 2581
rect 15 2439 25 2495
rect 81 2439 167 2495
rect 223 2439 309 2495
rect 365 2439 375 2495
rect 15 2353 375 2439
rect 15 2297 25 2353
rect 81 2297 167 2353
rect 223 2297 309 2353
rect 365 2297 375 2353
rect 15 2211 375 2297
rect 15 2155 25 2211
rect 81 2155 167 2211
rect 223 2155 309 2211
rect 365 2155 375 2211
rect 15 2069 375 2155
rect 15 2013 25 2069
rect 81 2013 167 2069
rect 223 2013 309 2069
rect 365 2013 375 2069
rect 15 1927 375 2013
rect 15 1871 25 1927
rect 81 1871 167 1927
rect 223 1871 309 1927
rect 365 1871 375 1927
rect 15 1785 375 1871
rect 15 1729 25 1785
rect 81 1729 167 1785
rect 223 1729 309 1785
rect 365 1729 375 1785
rect 15 1719 375 1729
rect 5523 2749 5883 2835
rect 5523 2693 5533 2749
rect 5589 2693 5675 2749
rect 5731 2693 5817 2749
rect 5873 2693 5883 2749
rect 5523 2607 5883 2693
rect 5523 2551 5533 2607
rect 5589 2551 5675 2607
rect 5731 2551 5817 2607
rect 5873 2551 5883 2607
rect 5523 2465 5883 2551
rect 5523 2409 5533 2465
rect 5589 2409 5675 2465
rect 5731 2409 5817 2465
rect 5873 2409 5883 2465
rect 5523 2323 5883 2409
rect 5523 2267 5533 2323
rect 5589 2267 5675 2323
rect 5731 2267 5817 2323
rect 5873 2267 5883 2323
rect 5523 2181 5883 2267
rect 5523 2125 5533 2181
rect 5589 2125 5675 2181
rect 5731 2125 5817 2181
rect 5873 2125 5883 2181
rect 5523 2039 5883 2125
rect 5523 1983 5533 2039
rect 5589 1983 5675 2039
rect 5731 1983 5817 2039
rect 5873 1983 5883 2039
rect 5523 1897 5883 1983
rect 5523 1841 5533 1897
rect 5589 1841 5675 1897
rect 5731 1841 5817 1897
rect 5873 1841 5883 1897
rect 5523 1755 5883 1841
rect 5523 1699 5533 1755
rect 5589 1699 5675 1755
rect 5731 1699 5817 1755
rect 5873 1699 5883 1755
rect 5523 1689 5883 1699
rect 550 1418 768 1428
rect 550 1362 560 1418
rect 616 1362 702 1418
rect 758 1362 768 1418
rect 550 1276 768 1362
rect 550 1220 560 1276
rect 616 1220 702 1276
rect 758 1220 768 1276
rect 550 1134 768 1220
rect 550 1078 560 1134
rect 616 1078 702 1134
rect 758 1078 768 1134
rect 550 992 768 1078
rect 550 936 560 992
rect 616 936 702 992
rect 758 936 768 992
rect 550 926 768 936
rect 1498 1418 1858 1428
rect 1498 1362 1508 1418
rect 1564 1362 1650 1418
rect 1706 1362 1792 1418
rect 1848 1362 1858 1418
rect 1498 1276 1858 1362
rect 1498 1220 1508 1276
rect 1564 1220 1650 1276
rect 1706 1220 1792 1276
rect 1848 1220 1858 1276
rect 1498 1134 1858 1220
rect 1498 1078 1508 1134
rect 1564 1078 1650 1134
rect 1706 1078 1792 1134
rect 1848 1078 1858 1134
rect 1498 992 1858 1078
rect 1498 936 1508 992
rect 1564 936 1650 992
rect 1706 936 1792 992
rect 1848 936 1858 992
rect 1498 926 1858 936
rect 2525 1418 2743 1428
rect 2525 1362 2535 1418
rect 2591 1362 2677 1418
rect 2733 1362 2743 1418
rect 2525 1276 2743 1362
rect 2525 1220 2535 1276
rect 2591 1220 2677 1276
rect 2733 1220 2743 1276
rect 2525 1134 2743 1220
rect 2525 1078 2535 1134
rect 2591 1078 2677 1134
rect 2733 1078 2743 1134
rect 2525 992 2743 1078
rect 2525 936 2535 992
rect 2591 936 2677 992
rect 2733 936 2743 992
rect 2525 926 2743 936
rect 3156 1418 3374 1428
rect 3156 1362 3166 1418
rect 3222 1362 3308 1418
rect 3364 1362 3374 1418
rect 3156 1276 3374 1362
rect 3156 1220 3166 1276
rect 3222 1220 3308 1276
rect 3364 1220 3374 1276
rect 3156 1134 3374 1220
rect 3156 1078 3166 1134
rect 3222 1078 3308 1134
rect 3364 1078 3374 1134
rect 3156 992 3374 1078
rect 3156 936 3166 992
rect 3222 936 3308 992
rect 3364 936 3374 992
rect 3156 926 3374 936
rect 4040 1418 4400 1428
rect 4040 1362 4050 1418
rect 4106 1362 4192 1418
rect 4248 1362 4334 1418
rect 4390 1362 4400 1418
rect 4040 1276 4400 1362
rect 4040 1220 4050 1276
rect 4106 1220 4192 1276
rect 4248 1220 4334 1276
rect 4390 1220 4400 1276
rect 4040 1134 4400 1220
rect 4040 1078 4050 1134
rect 4106 1078 4192 1134
rect 4248 1078 4334 1134
rect 4390 1078 4400 1134
rect 4040 992 4400 1078
rect 4040 936 4050 992
rect 4106 936 4192 992
rect 4248 936 4334 992
rect 4390 936 4400 992
rect 4040 926 4400 936
rect 5130 1418 5348 1428
rect 5130 1362 5140 1418
rect 5196 1362 5282 1418
rect 5338 1362 5348 1418
rect 5130 1276 5348 1362
rect 5130 1220 5140 1276
rect 5196 1220 5282 1276
rect 5338 1220 5348 1276
rect 5130 1134 5348 1220
rect 5130 1078 5140 1134
rect 5196 1078 5282 1134
rect 5338 1078 5348 1134
rect 5130 992 5348 1078
rect 5130 936 5140 992
rect 5196 936 5282 992
rect 5338 936 5348 992
rect 5130 926 5348 936
rect 568 787 2774 797
rect 568 731 578 787
rect 634 731 720 787
rect 776 731 862 787
rect 918 731 1004 787
rect 1060 731 1146 787
rect 1202 731 1288 787
rect 1344 731 1430 787
rect 1486 731 1572 787
rect 1628 731 1714 787
rect 1770 731 1856 787
rect 1912 731 1998 787
rect 2054 731 2140 787
rect 2196 731 2282 787
rect 2338 731 2424 787
rect 2480 731 2566 787
rect 2622 731 2708 787
rect 2764 731 2774 787
rect 568 645 2774 731
rect 568 589 578 645
rect 634 589 720 645
rect 776 589 862 645
rect 918 589 1004 645
rect 1060 589 1146 645
rect 1202 589 1288 645
rect 1344 589 1430 645
rect 1486 589 1572 645
rect 1628 589 1714 645
rect 1770 589 1856 645
rect 1912 589 1998 645
rect 2054 589 2140 645
rect 2196 589 2282 645
rect 2338 589 2424 645
rect 2480 589 2566 645
rect 2622 589 2708 645
rect 2764 589 2774 645
rect 568 579 2774 589
rect 3124 787 5330 797
rect 3124 731 3134 787
rect 3190 731 3276 787
rect 3332 731 3418 787
rect 3474 731 3560 787
rect 3616 731 3702 787
rect 3758 731 3844 787
rect 3900 731 3986 787
rect 4042 731 4128 787
rect 4184 731 4270 787
rect 4326 731 4412 787
rect 4468 731 4554 787
rect 4610 731 4696 787
rect 4752 731 4838 787
rect 4894 731 4980 787
rect 5036 731 5122 787
rect 5178 731 5264 787
rect 5320 731 5330 787
rect 3124 645 5330 731
rect 3124 589 3134 645
rect 3190 589 3276 645
rect 3332 589 3418 645
rect 3474 589 3560 645
rect 3616 589 3702 645
rect 3758 589 3844 645
rect 3900 589 3986 645
rect 4042 589 4128 645
rect 4184 589 4270 645
rect 4326 589 4412 645
rect 4468 589 4554 645
rect 4610 589 4696 645
rect 4752 589 4838 645
rect 4894 589 4980 645
rect 5036 589 5122 645
rect 5178 589 5264 645
rect 5320 589 5330 645
rect 3124 579 5330 589
use M1_NACTIVE_CDNS_40661956134345  M1_NACTIVE_CDNS_40661956134345_0
timestamp 1750858719
transform 1 0 2949 0 1 5716
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134345  M1_NACTIVE_CDNS_40661956134345_1
timestamp 1750858719
transform 1 0 2949 0 1 3848
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134346  M1_NACTIVE_CDNS_40661956134346_0
timestamp 1750858719
transform 1 0 5703 0 1 1545
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134346  M1_NACTIVE_CDNS_40661956134346_1
timestamp 1750858719
transform 1 0 195 0 1 1545
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134347  M1_NACTIVE_CDNS_40661956134347_0
timestamp 1750858719
transform 1 0 2949 0 1 4002
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134347  M1_NACTIVE_CDNS_40661956134347_1
timestamp 1750858719
transform 1 0 2949 0 1 4628
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134347  M1_NACTIVE_CDNS_40661956134347_2
timestamp 1750858719
transform 1 0 2949 0 1 5562
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134347  M1_NACTIVE_CDNS_40661956134347_3
timestamp 1750858719
transform 1 0 2949 0 1 4936
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134348  M1_NACTIVE_CDNS_40661956134348_0
timestamp 1750858719
transform 1 0 736 0 1 5252
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134348  M1_NACTIVE_CDNS_40661956134348_1
timestamp 1750858719
transform 1 0 5162 0 1 5252
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134348  M1_NACTIVE_CDNS_40661956134348_2
timestamp 1750858719
transform 1 0 736 0 1 4318
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134348  M1_NACTIVE_CDNS_40661956134348_3
timestamp 1750858719
transform 1 0 5162 0 1 4318
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134349  M1_NACTIVE_CDNS_40661956134349_0
timestamp 1750858719
transform 1 0 2949 0 1 4782
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134350  M1_NACTIVE_CDNS_40661956134350_0
timestamp 1750858719
transform 1 0 582 0 1 4782
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134350  M1_NACTIVE_CDNS_40661956134350_1
timestamp 1750858719
transform 1 0 5316 0 1 4782
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134358  M1_NACTIVE_CDNS_40661956134358_0
timestamp 1750858719
transform 1 0 195 0 1 7469
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134358  M1_NACTIVE_CDNS_40661956134358_1
timestamp 1750858719
transform 1 0 5703 0 1 7469
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134359  M1_NACTIVE_CDNS_40661956134359_0
timestamp 1750858719
transform 1 0 2949 0 1 195
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134359  M1_NACTIVE_CDNS_40661956134359_1
timestamp 1750858719
transform 1 0 2949 0 1 2895
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134359  M1_NACTIVE_CDNS_40661956134359_2
timestamp 1750858719
transform 1 0 2949 0 1 6669
box 0 0 1 1
use M1_NACTIVE_CDNS_40661956134359  M1_NACTIVE_CDNS_40661956134359_3
timestamp 1750858719
transform 1 0 2949 0 1 8269
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134344  M1_PACTIVE_CDNS_40661956134344_0
timestamp 1750858719
transform 1 0 195 0 1 4782
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134344  M1_PACTIVE_CDNS_40661956134344_1
timestamp 1750858719
transform 1 0 5703 0 1 4782
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134352  M1_PACTIVE_CDNS_40661956134352_0
timestamp 1750858719
transform 1 0 2949 0 1 611
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134352  M1_PACTIVE_CDNS_40661956134352_1
timestamp 1750858719
transform 1 0 2949 0 1 2479
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134353  M1_PACTIVE_CDNS_40661956134353_0
timestamp 1750858719
transform 1 0 5316 0 1 1545
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134353  M1_PACTIVE_CDNS_40661956134353_1
timestamp 1750858719
transform 1 0 582 0 1 1545
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134354  M1_PACTIVE_CDNS_40661956134354_0
timestamp 1750858719
transform 1 0 2949 0 1 765
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134354  M1_PACTIVE_CDNS_40661956134354_1
timestamp 1750858719
transform 1 0 2949 0 1 2325
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134354  M1_PACTIVE_CDNS_40661956134354_2
timestamp 1750858719
transform 1 0 2949 0 1 1391
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134354  M1_PACTIVE_CDNS_40661956134354_3
timestamp 1750858719
transform 1 0 2949 0 1 1699
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134355  M1_PACTIVE_CDNS_40661956134355_0
timestamp 1750858719
transform 1 0 5162 0 1 2015
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134355  M1_PACTIVE_CDNS_40661956134355_1
timestamp 1750858719
transform 1 0 5162 0 1 1081
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134355  M1_PACTIVE_CDNS_40661956134355_2
timestamp 1750858719
transform 1 0 736 0 1 1081
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134355  M1_PACTIVE_CDNS_40661956134355_3
timestamp 1750858719
transform 1 0 736 0 1 2015
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134356  M1_PACTIVE_CDNS_40661956134356_0
timestamp 1750858719
transform 1 0 2949 0 1 1545
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134357  M1_PACTIVE_CDNS_40661956134357_0
timestamp 1750858719
transform 1 0 2949 0 1 6132
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134357  M1_PACTIVE_CDNS_40661956134357_1
timestamp 1750858719
transform 1 0 2949 0 1 3432
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_0
timestamp 1750858719
transform 1 0 3265 0 1 2402
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_1
timestamp 1750858719
transform 1 0 2634 0 1 2402
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_0
timestamp 1750858719
transform 1 0 4220 0 1 1545
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_1
timestamp 1750858719
transform 1 0 1678 0 1 1545
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_2
timestamp 1750858719
transform 1 0 2690 0 1 4782
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_3
timestamp 1750858719
transform 1 0 1678 0 1 4782
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_4
timestamp 1750858719
transform 1 0 4220 0 1 4782
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_5
timestamp 1750858719
transform 1 0 3208 0 1 4782
box 0 0 1 1
use M2_M1_CDNS_40661956134343  M2_M1_CDNS_40661956134343_0
timestamp 1750858719
transform 1 0 2948 0 -1 7067
box 0 0 1 1
use M2_M1_CDNS_40661956134343  M2_M1_CDNS_40661956134343_1
timestamp 1750858719
transform 1 0 2948 0 1 7871
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_0
timestamp 1750858719
transform 1 0 4726 0 1 2012
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_1
timestamp 1750858719
transform 1 0 3714 0 1 2012
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_2
timestamp 1750858719
transform 1 0 4726 0 1 1078
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_3
timestamp 1750858719
transform 1 0 3714 0 1 1078
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_4
timestamp 1750858719
transform 1 0 3208 0 1 3925
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_5
timestamp 1750858719
transform 1 0 4220 0 1 3925
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_6
timestamp 1750858719
transform 1 0 4220 0 1 2402
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_7
timestamp 1750858719
transform 1 0 1678 0 1 3925
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_8
timestamp 1750858719
transform 1 0 2690 0 1 3925
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_9
timestamp 1750858719
transform 1 0 1678 0 1 2402
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_10
timestamp 1750858719
transform 1 0 1172 0 1 2012
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_11
timestamp 1750858719
transform 1 0 2184 0 1 2012
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_12
timestamp 1750858719
transform 1 0 1172 0 1 1078
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_13
timestamp 1750858719
transform 1 0 2184 0 1 1078
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_14
timestamp 1750858719
transform 1 0 1172 0 1 5249
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_15
timestamp 1750858719
transform 1 0 2184 0 1 5249
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_16
timestamp 1750858719
transform 1 0 1678 0 1 5639
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_17
timestamp 1750858719
transform 1 0 2690 0 1 5639
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_18
timestamp 1750858719
transform 1 0 4726 0 1 5249
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_19
timestamp 1750858719
transform 1 0 3714 0 1 5249
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_20
timestamp 1750858719
transform 1 0 3208 0 1 5639
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_21
timestamp 1750858719
transform 1 0 4220 0 1 5639
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_22
timestamp 1750858719
transform 1 0 1172 0 1 4315
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_23
timestamp 1750858719
transform 1 0 2184 0 1 4315
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_24
timestamp 1750858719
transform 1 0 4726 0 1 4315
box 0 0 1 1
use M2_M1_CDNS_40661956134351  M2_M1_CDNS_40661956134351_25
timestamp 1750858719
transform 1 0 3714 0 1 4315
box 0 0 1 1
use M2_M1_CDNS_40661956134360  M2_M1_CDNS_40661956134360_0
timestamp 1750858719
transform 1 0 3263 0 1 1545
box 0 0 1 1
use M2_M1_CDNS_40661956134360  M2_M1_CDNS_40661956134360_1
timestamp 1750858719
transform 1 0 2632 0 1 1545
box 0 0 1 1
use M2_M1_CDNS_40661956134361  M2_M1_CDNS_40661956134361_0
timestamp 1750858719
transform 1 0 5239 0 1 1012
box 0 0 1 1
use M2_M1_CDNS_40661956134361  M2_M1_CDNS_40661956134361_1
timestamp 1750858719
transform 1 0 659 0 1 1012
box 0 0 1 1
use M2_M1_CDNS_40661956134361  M2_M1_CDNS_40661956134361_2
timestamp 1750858719
transform 1 0 659 0 1 5304
box 0 0 1 1
use M2_M1_CDNS_40661956134361  M2_M1_CDNS_40661956134361_3
timestamp 1750858719
transform 1 0 5239 0 1 5304
box 0 0 1 1
use M2_M1_CDNS_40661956134363  M2_M1_CDNS_40661956134363_0
timestamp 1750858719
transform 1 0 195 0 1 4099
box 0 0 1 1
use M2_M1_CDNS_40661956134364  M2_M1_CDNS_40661956134364_0
timestamp 1750858719
transform 1 0 5703 0 1 2359
box 0 0 1 1
use M2_M1_CDNS_40661956134364  M2_M1_CDNS_40661956134364_1
timestamp 1750858719
transform 1 0 5703 0 1 3959
box 0 0 1 1
use M2_M1_CDNS_40661956134365  M2_M1_CDNS_40661956134365_0
timestamp 1750858719
transform 1 0 195 0 1 2255
box 0 0 1 1
use M2_M1_CDNS_40661956134370  M2_M1_CDNS_40661956134370_0
timestamp 1750858719
transform 1 0 1518 0 1 8269
box 0 0 1 1
use M2_M1_CDNS_40661956134370  M2_M1_CDNS_40661956134370_1
timestamp 1750858719
transform 1 0 4380 0 1 8269
box 0 0 1 1
use M2_M1_CDNS_40661956134371  M2_M1_CDNS_40661956134371_0
timestamp 1750858719
transform 0 1 195 -1 0 7469
box 0 0 1 1
use M2_M1_CDNS_40661956134371  M2_M1_CDNS_40661956134371_1
timestamp 1750858719
transform 0 1 5703 -1 0 7469
box 0 0 1 1
use M2_M1_CDNS_40661956134374  M2_M1_CDNS_40661956134374_0
timestamp 1750858719
transform 1 0 4137 0 1 688
box 0 0 1 1
use M2_M1_CDNS_40661956134374  M2_M1_CDNS_40661956134374_1
timestamp 1750858719
transform 1 0 1761 0 1 688
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_0
timestamp 1750858719
transform 1 0 5703 0 1 2366
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_1
timestamp 1750858719
transform 1 0 195 0 1 7168
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_2
timestamp 1750858719
transform 1 0 5703 0 1 7168
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_3
timestamp 1750858719
transform 1 0 5703 0 1 3959
box 0 0 1 1
use M3_M2_CDNS_40661956134362  M3_M2_CDNS_40661956134362_0
timestamp 1750858719
transform 1 0 4220 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134362  M3_M2_CDNS_40661956134362_1
timestamp 1750858719
transform 1 0 1678 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134366  M3_M2_CDNS_40661956134366_0
timestamp 1750858719
transform 1 0 2690 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134366  M3_M2_CDNS_40661956134366_1
timestamp 1750858719
transform 1 0 1678 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134366  M3_M2_CDNS_40661956134366_2
timestamp 1750858719
transform 1 0 3208 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134366  M3_M2_CDNS_40661956134366_3
timestamp 1750858719
transform 1 0 4220 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134367  M3_M2_CDNS_40661956134367_0
timestamp 1750858719
transform 1 0 195 0 1 2254
box 0 0 1 1
use M3_M2_CDNS_40661956134367  M3_M2_CDNS_40661956134367_1
timestamp 1750858719
transform 1 0 195 0 1 4099
box 0 0 1 1
use M3_M2_CDNS_40661956134368  M3_M2_CDNS_40661956134368_0
timestamp 1750858719
transform 1 0 3265 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134368  M3_M2_CDNS_40661956134368_1
timestamp 1750858719
transform 1 0 5239 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134368  M3_M2_CDNS_40661956134368_2
timestamp 1750858719
transform 1 0 2634 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134368  M3_M2_CDNS_40661956134368_3
timestamp 1750858719
transform 1 0 659 0 1 1177
box 0 0 1 1
use M3_M2_CDNS_40661956134369  M3_M2_CDNS_40661956134369_0
timestamp 1750858719
transform 1 0 1260 0 1 8269
box 0 0 1 1
use M3_M2_CDNS_40661956134369  M3_M2_CDNS_40661956134369_1
timestamp 1750858719
transform 1 0 4638 0 1 8269
box 0 0 1 1
use M3_M2_CDNS_40661956134372  M3_M2_CDNS_40661956134372_0
timestamp 1750858719
transform 1 0 659 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134372  M3_M2_CDNS_40661956134372_1
timestamp 1750858719
transform 1 0 5239 0 1 5305
box 0 0 1 1
use M3_M2_CDNS_40661956134373  M3_M2_CDNS_40661956134373_0
timestamp 1750858719
transform 1 0 4227 0 1 688
box 0 0 1 1
use M3_M2_CDNS_40661956134373  M3_M2_CDNS_40661956134373_1
timestamp 1750858719
transform 1 0 1671 0 1 688
box 0 0 1 1
use np_6p0_CDNS_4066195613426  np_6p0_CDNS_4066195613426_0
timestamp 1750858719
transform 0 1 949 -1 0 2112
box 0 0 1 1
use np_6p0_CDNS_4066195613426  np_6p0_CDNS_4066195613426_1
timestamp 1750858719
transform 0 1 949 -1 0 1178
box 0 0 1 1
use pn_6p0_CDNS_4066195613427  pn_6p0_CDNS_4066195613427_0
timestamp 1750858719
transform 0 1 949 -1 0 4415
box 0 0 1 1
use pn_6p0_CDNS_4066195613427  pn_6p0_CDNS_4066195613427_1
timestamp 1750858719
transform 0 1 949 -1 0 5349
box 0 0 1 1
use ppolyf_u_CDNS_4066195613425  ppolyf_u_CDNS_4066195613425_0
timestamp 1750858719
transform 0 1 1769 -1 0 7851
box 0 0 1 1
use ppolyf_u_CDNS_4066195613425  ppolyf_u_CDNS_4066195613425_1
timestamp 1750858719
transform 0 1 2389 -1 0 7851
box 0 0 1 1
use ppolyf_u_CDNS_4066195613425  ppolyf_u_CDNS_4066195613425_2
timestamp 1750858719
transform 0 1 3629 -1 0 7851
box 0 0 1 1
use ppolyf_u_CDNS_4066195613425  ppolyf_u_CDNS_4066195613425_3
timestamp 1750858719
transform 0 1 3009 -1 0 7851
box 0 0 1 1
<< labels >>
rlabel metal2 s 2965 6784 2965 6784 4 IP_IN
port 1 nsew
rlabel metal2 s 2965 7877 2965 7877 4 PAD
port 2 nsew
rlabel metal1 s 494 8257 494 8257 4 DVDD
port 3 nsew
rlabel metal1 s 494 6132 494 6132 4 DVSS
port 4 nsew
<< properties >>
string GDS_END 879400
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 868170
string path 123.725 79.725 -5.125 79.725 
<< end >>
