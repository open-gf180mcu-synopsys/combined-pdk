magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 1800 1660
<< nmos >>
rect 200 210 260 380
rect 400 210 460 380
rect 540 210 600 380
rect 710 210 770 380
rect 850 210 910 380
rect 1050 210 1110 380
rect 1370 210 1430 380
rect 1540 210 1600 380
<< pmos >>
rect 200 1110 260 1450
rect 370 1110 430 1450
rect 540 1110 600 1450
rect 710 1110 770 1450
rect 880 1110 940 1450
rect 1050 1110 1110 1450
rect 1370 1110 1430 1450
rect 1540 1110 1600 1450
<< ndiff >>
rect 100 318 200 380
rect 100 272 122 318
rect 168 272 200 318
rect 100 210 200 272
rect 260 318 400 380
rect 260 272 307 318
rect 353 272 400 318
rect 260 210 400 272
rect 460 210 540 380
rect 600 318 710 380
rect 600 272 632 318
rect 678 272 710 318
rect 600 210 710 272
rect 770 210 850 380
rect 910 318 1050 380
rect 910 272 957 318
rect 1003 272 1050 318
rect 910 210 1050 272
rect 1110 318 1210 380
rect 1110 272 1142 318
rect 1188 272 1210 318
rect 1110 210 1210 272
rect 1270 318 1370 380
rect 1270 272 1292 318
rect 1338 272 1370 318
rect 1270 210 1370 272
rect 1430 318 1540 380
rect 1430 272 1462 318
rect 1508 272 1540 318
rect 1430 210 1540 272
rect 1600 318 1700 380
rect 1600 272 1632 318
rect 1678 272 1700 318
rect 1600 210 1700 272
<< pdiff >>
rect 100 1397 200 1450
rect 100 1163 122 1397
rect 168 1163 200 1397
rect 100 1110 200 1163
rect 260 1430 370 1450
rect 260 1290 292 1430
rect 338 1290 370 1430
rect 260 1110 370 1290
rect 430 1110 540 1450
rect 600 1397 710 1450
rect 600 1163 632 1397
rect 678 1163 710 1397
rect 600 1110 710 1163
rect 770 1110 880 1450
rect 940 1397 1050 1450
rect 940 1163 972 1397
rect 1018 1163 1050 1397
rect 940 1110 1050 1163
rect 1110 1397 1210 1450
rect 1110 1163 1142 1397
rect 1188 1163 1210 1397
rect 1110 1110 1210 1163
rect 1270 1397 1370 1450
rect 1270 1163 1292 1397
rect 1338 1163 1370 1397
rect 1270 1110 1370 1163
rect 1430 1397 1540 1450
rect 1430 1163 1462 1397
rect 1508 1163 1540 1397
rect 1430 1110 1540 1163
rect 1600 1397 1700 1450
rect 1600 1163 1632 1397
rect 1678 1163 1700 1397
rect 1600 1110 1700 1163
<< ndiffc >>
rect 122 272 168 318
rect 307 272 353 318
rect 632 272 678 318
rect 957 272 1003 318
rect 1142 272 1188 318
rect 1292 272 1338 318
rect 1462 272 1508 318
rect 1632 272 1678 318
<< pdiffc >>
rect 122 1163 168 1397
rect 292 1290 338 1430
rect 632 1163 678 1397
rect 972 1163 1018 1397
rect 1142 1163 1188 1397
rect 1292 1163 1338 1397
rect 1462 1163 1508 1397
rect 1632 1163 1678 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1030 118 1180 140
rect 1030 72 1082 118
rect 1128 72 1180 118
rect 1030 50 1180 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 310 1588 460 1610
rect 310 1542 362 1588
rect 408 1542 460 1588
rect 310 1520 460 1542
rect 540 1588 690 1610
rect 540 1542 592 1588
rect 638 1542 690 1588
rect 540 1520 690 1542
rect 780 1588 930 1610
rect 780 1542 832 1588
rect 878 1542 930 1588
rect 780 1520 930 1542
rect 1030 1588 1180 1610
rect 1030 1542 1082 1588
rect 1128 1542 1180 1588
rect 1030 1520 1180 1542
rect 1270 1588 1420 1610
rect 1270 1542 1322 1588
rect 1368 1542 1420 1588
rect 1270 1520 1420 1542
rect 1510 1588 1660 1610
rect 1510 1542 1562 1588
rect 1608 1542 1660 1588
rect 1510 1520 1660 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 592 72 638 118
rect 832 72 878 118
rect 1082 72 1128 118
rect 1312 72 1358 118
rect 1552 72 1598 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 362 1542 408 1588
rect 592 1542 638 1588
rect 832 1542 878 1588
rect 1082 1542 1128 1588
rect 1322 1542 1368 1588
rect 1562 1542 1608 1588
<< polysilicon >>
rect 200 1450 260 1500
rect 370 1450 430 1500
rect 540 1450 600 1500
rect 710 1450 770 1500
rect 880 1450 940 1500
rect 1050 1450 1110 1500
rect 1370 1450 1430 1500
rect 1540 1450 1600 1500
rect 200 930 260 1110
rect 370 930 430 1110
rect 540 1040 600 1110
rect 520 1013 620 1040
rect 520 967 547 1013
rect 593 967 620 1013
rect 520 940 620 967
rect 710 930 770 1110
rect 200 903 320 930
rect 200 857 237 903
rect 283 857 320 903
rect 200 830 320 857
rect 370 903 470 930
rect 370 857 397 903
rect 443 857 470 903
rect 370 830 470 857
rect 690 903 790 930
rect 690 857 717 903
rect 763 857 790 903
rect 690 830 790 857
rect 200 380 260 830
rect 370 470 430 830
rect 710 720 770 830
rect 540 660 770 720
rect 880 800 940 1110
rect 1050 930 1110 1110
rect 1040 903 1140 930
rect 1040 857 1067 903
rect 1113 857 1140 903
rect 1040 830 1140 857
rect 880 773 1000 800
rect 880 727 927 773
rect 973 727 1000 773
rect 880 700 1000 727
rect 370 430 460 470
rect 400 380 460 430
rect 540 380 600 660
rect 690 583 790 610
rect 690 537 717 583
rect 763 537 790 583
rect 690 510 790 537
rect 710 380 770 510
rect 880 470 940 700
rect 850 430 940 470
rect 850 380 910 430
rect 1050 380 1110 830
rect 1370 800 1430 1110
rect 1540 930 1600 1110
rect 1480 903 1600 930
rect 1480 857 1507 903
rect 1553 857 1600 903
rect 1480 830 1600 857
rect 1350 778 1440 800
rect 1350 732 1372 778
rect 1418 732 1440 778
rect 1350 710 1440 732
rect 1370 380 1430 710
rect 1540 380 1600 830
rect 200 160 260 210
rect 400 160 460 210
rect 540 160 600 210
rect 710 160 770 210
rect 850 160 910 210
rect 1050 160 1110 210
rect 1370 160 1430 210
rect 1540 160 1600 210
<< polycontact >>
rect 547 967 593 1013
rect 237 857 283 903
rect 397 857 443 903
rect 717 857 763 903
rect 1067 857 1113 903
rect 927 727 973 773
rect 717 537 763 583
rect 1507 857 1553 903
rect 1372 732 1418 778
<< metal1 >>
rect 0 1588 1800 1660
rect 0 1542 112 1588
rect 158 1542 362 1588
rect 408 1542 592 1588
rect 638 1542 832 1588
rect 878 1542 1082 1588
rect 1128 1542 1322 1588
rect 1368 1542 1562 1588
rect 1608 1542 1800 1588
rect 0 1520 1800 1542
rect 120 1397 170 1450
rect 120 1163 122 1397
rect 168 1163 170 1397
rect 290 1430 340 1520
rect 290 1290 292 1430
rect 338 1290 340 1430
rect 290 1270 340 1290
rect 630 1397 680 1450
rect 120 790 170 1163
rect 630 1163 632 1397
rect 678 1163 680 1397
rect 630 1160 680 1163
rect 230 1110 680 1160
rect 970 1397 1020 1520
rect 970 1163 972 1397
rect 1018 1163 1020 1397
rect 970 1110 1020 1163
rect 1140 1397 1190 1450
rect 1140 1163 1142 1397
rect 1188 1163 1190 1397
rect 1140 1120 1190 1163
rect 1290 1397 1340 1450
rect 1290 1163 1292 1397
rect 1338 1163 1340 1397
rect 230 910 280 1110
rect 1140 1070 1240 1120
rect 520 1013 620 1020
rect 520 967 547 1013
rect 593 967 620 1013
rect 520 960 620 967
rect 220 903 310 910
rect 220 857 237 903
rect 283 857 310 903
rect 220 850 310 857
rect 370 906 470 910
rect 370 854 394 906
rect 446 854 470 906
rect 370 850 470 854
rect 100 780 170 790
rect 70 776 170 780
rect 70 724 94 776
rect 146 724 170 776
rect 70 720 170 724
rect 90 710 170 720
rect 120 318 170 710
rect 230 480 280 850
rect 540 590 600 960
rect 690 906 790 910
rect 690 854 714 906
rect 766 854 790 906
rect 690 850 790 854
rect 1040 906 1140 910
rect 1040 854 1064 906
rect 1116 854 1140 906
rect 1040 850 1140 854
rect 900 776 1000 780
rect 900 724 924 776
rect 976 724 1000 776
rect 900 720 1000 724
rect 1190 590 1240 1070
rect 1290 1080 1340 1163
rect 1460 1397 1510 1520
rect 1460 1163 1462 1397
rect 1508 1163 1510 1397
rect 1460 1110 1510 1163
rect 1630 1397 1680 1450
rect 1630 1163 1632 1397
rect 1678 1163 1680 1397
rect 1290 1040 1370 1080
rect 1630 1050 1680 1163
rect 1630 1040 1710 1050
rect 1290 1036 1390 1040
rect 1290 984 1314 1036
rect 1366 1030 1390 1036
rect 1630 1036 1730 1040
rect 1366 984 1560 1030
rect 1290 980 1560 984
rect 1290 970 1370 980
rect 1500 903 1560 980
rect 1500 857 1507 903
rect 1553 857 1560 903
rect 1350 778 1450 780
rect 1350 732 1372 778
rect 1418 776 1450 778
rect 1350 724 1374 732
rect 1426 724 1450 776
rect 1350 720 1450 724
rect 540 583 1240 590
rect 540 537 717 583
rect 763 537 1240 583
rect 540 530 1240 537
rect 230 430 680 480
rect 1190 460 1240 530
rect 1500 480 1560 857
rect 120 272 122 318
rect 168 272 170 318
rect 120 210 170 272
rect 290 318 370 380
rect 290 272 307 318
rect 353 272 370 318
rect 290 140 370 272
rect 630 318 680 430
rect 1140 410 1240 460
rect 1290 430 1560 480
rect 1630 984 1654 1036
rect 1706 984 1730 1036
rect 1630 980 1730 984
rect 1630 970 1710 980
rect 630 272 632 318
rect 678 272 680 318
rect 630 210 680 272
rect 940 318 1020 380
rect 940 272 957 318
rect 1003 272 1020 318
rect 940 140 1020 272
rect 1140 318 1190 410
rect 1140 272 1142 318
rect 1188 272 1190 318
rect 1140 210 1190 272
rect 1290 318 1340 430
rect 1290 272 1292 318
rect 1338 272 1340 318
rect 1290 210 1340 272
rect 1460 318 1510 380
rect 1460 272 1462 318
rect 1508 272 1510 318
rect 1460 140 1510 272
rect 1630 318 1680 970
rect 1630 272 1632 318
rect 1678 272 1680 318
rect 1630 210 1680 272
rect 0 118 1800 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 592 118
rect 638 72 832 118
rect 878 72 1082 118
rect 1128 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1800 118
rect 0 0 1800 72
<< via1 >>
rect 394 903 446 906
rect 394 857 397 903
rect 397 857 443 903
rect 443 857 446 903
rect 394 854 446 857
rect 94 724 146 776
rect 714 903 766 906
rect 714 857 717 903
rect 717 857 763 903
rect 763 857 766 903
rect 714 854 766 857
rect 1064 903 1116 906
rect 1064 857 1067 903
rect 1067 857 1113 903
rect 1113 857 1116 903
rect 1064 854 1116 857
rect 924 773 976 776
rect 924 727 927 773
rect 927 727 973 773
rect 973 727 976 773
rect 924 724 976 727
rect 1314 984 1366 1036
rect 1374 732 1418 776
rect 1418 732 1426 776
rect 1374 724 1426 732
rect 1654 984 1706 1036
<< metal2 >>
rect 1300 1040 1380 1050
rect 1640 1040 1720 1050
rect 1290 1036 1390 1040
rect 1290 984 1314 1036
rect 1366 984 1390 1036
rect 1290 980 1390 984
rect 1630 1036 1730 1040
rect 1630 984 1654 1036
rect 1706 984 1730 1036
rect 1630 980 1730 984
rect 1300 970 1380 980
rect 1640 970 1720 980
rect 370 906 470 920
rect 700 910 780 920
rect 1040 910 1140 920
rect 370 854 394 906
rect 446 854 470 906
rect 370 840 470 854
rect 690 906 1140 910
rect 690 854 714 906
rect 766 854 1064 906
rect 1116 854 1140 906
rect 690 850 1140 854
rect 700 840 780 850
rect 1040 840 1140 850
rect 70 780 170 790
rect 910 780 990 790
rect 1350 780 1450 790
rect 70 776 1450 780
rect 70 724 94 776
rect 146 724 924 776
rect 976 724 1374 776
rect 1426 724 1450 776
rect 70 720 1450 724
rect 70 710 170 720
rect 910 710 990 720
rect 1350 710 1450 720
<< labels >>
rlabel via1 s 394 854 446 906 4 D
port 1 nsew signal input
rlabel via1 s 1654 984 1706 1036 4 Q
port 2 nsew signal output
rlabel via1 s 1064 854 1116 906 4 CLK
port 3 nsew clock input
rlabel metal1 s 290 1270 340 1660 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 0 370 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 714 854 766 906 1 CLK
port 3 nsew clock input
rlabel metal1 s 690 850 790 910 1 CLK
port 3 nsew clock input
rlabel metal1 s 1040 850 1140 910 1 CLK
port 3 nsew clock input
rlabel metal2 s 700 840 780 920 1 CLK
port 3 nsew clock input
rlabel metal2 s 690 850 1140 910 1 CLK
port 3 nsew clock input
rlabel metal2 s 1040 840 1140 920 1 CLK
port 3 nsew clock input
rlabel metal1 s 970 1110 1020 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1460 1110 1510 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1520 1800 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 940 0 1020 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1460 0 1510 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1800 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 370 850 470 910 1 D
port 1 nsew signal input
rlabel metal2 s 370 840 470 920 1 D
port 1 nsew signal input
rlabel metal1 s 1630 210 1680 1450 1 Q
port 2 nsew signal output
rlabel metal1 s 1630 970 1710 1050 1 Q
port 2 nsew signal output
rlabel metal1 s 1630 980 1730 1040 1 Q
port 2 nsew signal output
rlabel metal2 s 1640 970 1720 1050 1 Q
port 2 nsew signal output
rlabel metal2 s 1630 980 1730 1040 1 Q
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1800 1660
string GDS_END 388160
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 375224
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
