magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -1030 29053 21660 29790
<< mvpmos >>
rect -754 29194 -281 29649
rect -135 29194 338 29649
rect 484 29194 957 29649
rect 1103 29194 1576 29649
rect 1722 29194 2195 29649
rect 2341 29194 2814 29649
rect 2960 29194 3433 29649
rect 3579 29194 4052 29649
rect 4198 29194 4671 29649
rect 4817 29194 5290 29649
rect 5436 29194 5909 29649
rect 6055 29194 6528 29649
rect 6674 29194 7147 29649
rect 7293 29194 7766 29649
rect 7912 29194 8385 29649
rect 8531 29194 9004 29649
rect 9150 29194 9623 29649
rect 9769 29194 10242 29649
rect 10388 29194 10861 29649
rect 11007 29194 11480 29649
rect 11626 29194 12099 29649
rect 12245 29194 12718 29649
rect 12864 29194 13337 29649
rect 13483 29194 13956 29649
rect 14102 29194 14575 29649
rect 14721 29194 15194 29649
rect 15340 29194 15813 29649
rect 15959 29194 16432 29649
rect 16578 29194 17051 29649
rect 17197 29194 17670 29649
rect 17816 29194 18289 29649
rect 18435 29194 18908 29649
rect 19054 29194 19527 29649
rect 19673 29194 20146 29649
rect 20292 29194 20765 29649
rect 20911 29194 21384 29649
<< mvpdiff >>
rect -894 29604 -754 29649
rect -894 29558 -850 29604
rect -804 29558 -754 29604
rect -894 29286 -754 29558
rect -894 29240 -850 29286
rect -804 29240 -754 29286
rect -894 29194 -754 29240
rect -281 29604 -135 29649
rect -281 29558 -231 29604
rect -185 29558 -135 29604
rect -281 29286 -135 29558
rect -281 29240 -231 29286
rect -185 29240 -135 29286
rect -281 29194 -135 29240
rect 338 29604 484 29649
rect 338 29558 388 29604
rect 434 29558 484 29604
rect 338 29286 484 29558
rect 338 29240 388 29286
rect 434 29240 484 29286
rect 338 29194 484 29240
rect 957 29604 1103 29649
rect 957 29558 1007 29604
rect 1053 29558 1103 29604
rect 957 29286 1103 29558
rect 957 29240 1007 29286
rect 1053 29240 1103 29286
rect 957 29194 1103 29240
rect 1576 29604 1722 29649
rect 1576 29558 1626 29604
rect 1672 29558 1722 29604
rect 1576 29286 1722 29558
rect 1576 29240 1626 29286
rect 1672 29240 1722 29286
rect 1576 29194 1722 29240
rect 2195 29604 2341 29649
rect 2195 29558 2245 29604
rect 2291 29558 2341 29604
rect 2195 29286 2341 29558
rect 2195 29240 2245 29286
rect 2291 29240 2341 29286
rect 2195 29194 2341 29240
rect 2814 29604 2960 29649
rect 2814 29558 2864 29604
rect 2910 29558 2960 29604
rect 2814 29286 2960 29558
rect 2814 29240 2864 29286
rect 2910 29240 2960 29286
rect 2814 29194 2960 29240
rect 3433 29604 3579 29649
rect 3433 29558 3483 29604
rect 3529 29558 3579 29604
rect 3433 29286 3579 29558
rect 3433 29240 3483 29286
rect 3529 29240 3579 29286
rect 3433 29194 3579 29240
rect 4052 29604 4198 29649
rect 4052 29558 4102 29604
rect 4148 29558 4198 29604
rect 4052 29286 4198 29558
rect 4052 29240 4102 29286
rect 4148 29240 4198 29286
rect 4052 29194 4198 29240
rect 4671 29604 4817 29649
rect 4671 29558 4721 29604
rect 4767 29558 4817 29604
rect 4671 29286 4817 29558
rect 4671 29240 4721 29286
rect 4767 29240 4817 29286
rect 4671 29194 4817 29240
rect 5290 29604 5436 29649
rect 5290 29558 5340 29604
rect 5386 29558 5436 29604
rect 5290 29286 5436 29558
rect 5290 29240 5340 29286
rect 5386 29240 5436 29286
rect 5290 29194 5436 29240
rect 5909 29604 6055 29649
rect 5909 29558 5959 29604
rect 6005 29558 6055 29604
rect 5909 29286 6055 29558
rect 5909 29240 5959 29286
rect 6005 29240 6055 29286
rect 5909 29194 6055 29240
rect 6528 29604 6674 29649
rect 6528 29558 6578 29604
rect 6624 29558 6674 29604
rect 6528 29286 6674 29558
rect 6528 29240 6578 29286
rect 6624 29240 6674 29286
rect 6528 29194 6674 29240
rect 7147 29604 7293 29649
rect 7147 29558 7197 29604
rect 7243 29558 7293 29604
rect 7147 29286 7293 29558
rect 7147 29240 7197 29286
rect 7243 29240 7293 29286
rect 7147 29194 7293 29240
rect 7766 29604 7912 29649
rect 7766 29558 7816 29604
rect 7862 29558 7912 29604
rect 7766 29286 7912 29558
rect 7766 29240 7816 29286
rect 7862 29240 7912 29286
rect 7766 29194 7912 29240
rect 8385 29604 8531 29649
rect 8385 29558 8435 29604
rect 8481 29558 8531 29604
rect 8385 29286 8531 29558
rect 8385 29240 8435 29286
rect 8481 29240 8531 29286
rect 8385 29194 8531 29240
rect 9004 29604 9150 29649
rect 9004 29558 9054 29604
rect 9100 29558 9150 29604
rect 9004 29286 9150 29558
rect 9004 29240 9054 29286
rect 9100 29240 9150 29286
rect 9004 29194 9150 29240
rect 9623 29604 9769 29649
rect 9623 29558 9673 29604
rect 9719 29558 9769 29604
rect 9623 29286 9769 29558
rect 9623 29240 9673 29286
rect 9719 29240 9769 29286
rect 9623 29194 9769 29240
rect 10242 29604 10388 29649
rect 10242 29558 10292 29604
rect 10338 29558 10388 29604
rect 10242 29286 10388 29558
rect 10242 29240 10292 29286
rect 10338 29240 10388 29286
rect 10242 29194 10388 29240
rect 10861 29604 11007 29649
rect 10861 29558 10911 29604
rect 10957 29558 11007 29604
rect 10861 29286 11007 29558
rect 10861 29240 10911 29286
rect 10957 29240 11007 29286
rect 10861 29194 11007 29240
rect 11480 29604 11626 29649
rect 11480 29558 11530 29604
rect 11576 29558 11626 29604
rect 11480 29286 11626 29558
rect 11480 29240 11530 29286
rect 11576 29240 11626 29286
rect 11480 29194 11626 29240
rect 12099 29604 12245 29649
rect 12099 29558 12149 29604
rect 12195 29558 12245 29604
rect 12099 29286 12245 29558
rect 12099 29240 12149 29286
rect 12195 29240 12245 29286
rect 12099 29194 12245 29240
rect 12718 29604 12864 29649
rect 12718 29558 12768 29604
rect 12814 29558 12864 29604
rect 12718 29286 12864 29558
rect 12718 29240 12768 29286
rect 12814 29240 12864 29286
rect 12718 29194 12864 29240
rect 13337 29604 13483 29649
rect 13337 29558 13387 29604
rect 13433 29558 13483 29604
rect 13337 29286 13483 29558
rect 13337 29240 13387 29286
rect 13433 29240 13483 29286
rect 13337 29194 13483 29240
rect 13956 29604 14102 29649
rect 13956 29558 14006 29604
rect 14052 29558 14102 29604
rect 13956 29286 14102 29558
rect 13956 29240 14006 29286
rect 14052 29240 14102 29286
rect 13956 29194 14102 29240
rect 14575 29604 14721 29649
rect 14575 29558 14625 29604
rect 14671 29558 14721 29604
rect 14575 29286 14721 29558
rect 14575 29240 14625 29286
rect 14671 29240 14721 29286
rect 14575 29194 14721 29240
rect 15194 29604 15340 29649
rect 15194 29558 15244 29604
rect 15290 29558 15340 29604
rect 15194 29286 15340 29558
rect 15194 29240 15244 29286
rect 15290 29240 15340 29286
rect 15194 29194 15340 29240
rect 15813 29604 15959 29649
rect 15813 29558 15863 29604
rect 15909 29558 15959 29604
rect 15813 29286 15959 29558
rect 15813 29240 15863 29286
rect 15909 29240 15959 29286
rect 15813 29194 15959 29240
rect 16432 29604 16578 29649
rect 16432 29558 16482 29604
rect 16528 29558 16578 29604
rect 16432 29286 16578 29558
rect 16432 29240 16482 29286
rect 16528 29240 16578 29286
rect 16432 29194 16578 29240
rect 17051 29604 17197 29649
rect 17051 29558 17101 29604
rect 17147 29558 17197 29604
rect 17051 29286 17197 29558
rect 17051 29240 17101 29286
rect 17147 29240 17197 29286
rect 17051 29194 17197 29240
rect 17670 29604 17816 29649
rect 17670 29558 17720 29604
rect 17766 29558 17816 29604
rect 17670 29286 17816 29558
rect 17670 29240 17720 29286
rect 17766 29240 17816 29286
rect 17670 29194 17816 29240
rect 18289 29604 18435 29649
rect 18289 29558 18339 29604
rect 18385 29558 18435 29604
rect 18289 29286 18435 29558
rect 18289 29240 18339 29286
rect 18385 29240 18435 29286
rect 18289 29194 18435 29240
rect 18908 29604 19054 29649
rect 18908 29558 18958 29604
rect 19004 29558 19054 29604
rect 18908 29286 19054 29558
rect 18908 29240 18958 29286
rect 19004 29240 19054 29286
rect 18908 29194 19054 29240
rect 19527 29604 19673 29649
rect 19527 29558 19577 29604
rect 19623 29558 19673 29604
rect 19527 29286 19673 29558
rect 19527 29240 19577 29286
rect 19623 29240 19673 29286
rect 19527 29194 19673 29240
rect 20146 29604 20292 29649
rect 20146 29558 20196 29604
rect 20242 29558 20292 29604
rect 20146 29286 20292 29558
rect 20146 29240 20196 29286
rect 20242 29240 20292 29286
rect 20146 29194 20292 29240
rect 20765 29604 20911 29649
rect 20765 29558 20815 29604
rect 20861 29558 20911 29604
rect 20765 29286 20911 29558
rect 20765 29240 20815 29286
rect 20861 29240 20911 29286
rect 20765 29194 20911 29240
rect 21384 29604 21524 29649
rect 21384 29558 21434 29604
rect 21480 29558 21524 29604
rect 21384 29286 21524 29558
rect 21384 29240 21434 29286
rect 21480 29240 21524 29286
rect 21384 29194 21524 29240
<< mvpdiffc >>
rect -850 29558 -804 29604
rect -850 29240 -804 29286
rect -231 29558 -185 29604
rect -231 29240 -185 29286
rect 388 29558 434 29604
rect 388 29240 434 29286
rect 1007 29558 1053 29604
rect 1007 29240 1053 29286
rect 1626 29558 1672 29604
rect 1626 29240 1672 29286
rect 2245 29558 2291 29604
rect 2245 29240 2291 29286
rect 2864 29558 2910 29604
rect 2864 29240 2910 29286
rect 3483 29558 3529 29604
rect 3483 29240 3529 29286
rect 4102 29558 4148 29604
rect 4102 29240 4148 29286
rect 4721 29558 4767 29604
rect 4721 29240 4767 29286
rect 5340 29558 5386 29604
rect 5340 29240 5386 29286
rect 5959 29558 6005 29604
rect 5959 29240 6005 29286
rect 6578 29558 6624 29604
rect 6578 29240 6624 29286
rect 7197 29558 7243 29604
rect 7197 29240 7243 29286
rect 7816 29558 7862 29604
rect 7816 29240 7862 29286
rect 8435 29558 8481 29604
rect 8435 29240 8481 29286
rect 9054 29558 9100 29604
rect 9054 29240 9100 29286
rect 9673 29558 9719 29604
rect 9673 29240 9719 29286
rect 10292 29558 10338 29604
rect 10292 29240 10338 29286
rect 10911 29558 10957 29604
rect 10911 29240 10957 29286
rect 11530 29558 11576 29604
rect 11530 29240 11576 29286
rect 12149 29558 12195 29604
rect 12149 29240 12195 29286
rect 12768 29558 12814 29604
rect 12768 29240 12814 29286
rect 13387 29558 13433 29604
rect 13387 29240 13433 29286
rect 14006 29558 14052 29604
rect 14006 29240 14052 29286
rect 14625 29558 14671 29604
rect 14625 29240 14671 29286
rect 15244 29558 15290 29604
rect 15244 29240 15290 29286
rect 15863 29558 15909 29604
rect 15863 29240 15909 29286
rect 16482 29558 16528 29604
rect 16482 29240 16528 29286
rect 17101 29558 17147 29604
rect 17101 29240 17147 29286
rect 17720 29558 17766 29604
rect 17720 29240 17766 29286
rect 18339 29558 18385 29604
rect 18339 29240 18385 29286
rect 18958 29558 19004 29604
rect 18958 29240 19004 29286
rect 19577 29558 19623 29604
rect 19577 29240 19623 29286
rect 20196 29558 20242 29604
rect 20196 29240 20242 29286
rect 20815 29558 20861 29604
rect 20815 29240 20861 29286
rect 21434 29558 21480 29604
rect 21434 29240 21480 29286
<< polysilicon >>
rect -754 29803 -281 29858
rect -754 29757 -701 29803
rect -655 29757 -380 29803
rect -334 29757 -281 29803
rect -754 29649 -281 29757
rect -135 29803 338 29858
rect -135 29757 -82 29803
rect -36 29757 239 29803
rect 285 29757 338 29803
rect -135 29649 338 29757
rect 484 29803 957 29858
rect 484 29757 537 29803
rect 583 29757 858 29803
rect 904 29757 957 29803
rect 484 29649 957 29757
rect 1103 29803 1576 29858
rect 1103 29757 1156 29803
rect 1202 29757 1477 29803
rect 1523 29757 1576 29803
rect 1103 29649 1576 29757
rect 1722 29803 2195 29858
rect 1722 29757 1775 29803
rect 1821 29757 2096 29803
rect 2142 29757 2195 29803
rect 1722 29649 2195 29757
rect 2341 29803 2814 29858
rect 2341 29757 2394 29803
rect 2440 29757 2715 29803
rect 2761 29757 2814 29803
rect 2341 29649 2814 29757
rect 2960 29803 3433 29858
rect 2960 29757 3013 29803
rect 3059 29757 3334 29803
rect 3380 29757 3433 29803
rect 2960 29649 3433 29757
rect 3579 29803 4052 29858
rect 3579 29757 3632 29803
rect 3678 29757 3953 29803
rect 3999 29757 4052 29803
rect 3579 29649 4052 29757
rect 4198 29803 4671 29858
rect 4198 29757 4251 29803
rect 4297 29757 4572 29803
rect 4618 29757 4671 29803
rect 4198 29649 4671 29757
rect 4817 29803 5290 29858
rect 4817 29757 4870 29803
rect 4916 29757 5191 29803
rect 5237 29757 5290 29803
rect 4817 29649 5290 29757
rect 5436 29803 5909 29858
rect 5436 29757 5489 29803
rect 5535 29757 5810 29803
rect 5856 29757 5909 29803
rect 5436 29649 5909 29757
rect 6055 29803 6528 29858
rect 6055 29757 6108 29803
rect 6154 29757 6429 29803
rect 6475 29757 6528 29803
rect 6055 29649 6528 29757
rect 6674 29803 7147 29858
rect 6674 29757 6727 29803
rect 6773 29757 7048 29803
rect 7094 29757 7147 29803
rect 6674 29649 7147 29757
rect 7293 29803 7766 29858
rect 7293 29757 7346 29803
rect 7392 29757 7667 29803
rect 7713 29757 7766 29803
rect 7293 29649 7766 29757
rect 7912 29803 8385 29858
rect 7912 29757 7965 29803
rect 8011 29757 8286 29803
rect 8332 29757 8385 29803
rect 7912 29649 8385 29757
rect 8531 29803 9004 29858
rect 8531 29757 8584 29803
rect 8630 29757 8905 29803
rect 8951 29757 9004 29803
rect 8531 29649 9004 29757
rect 9150 29803 9623 29858
rect 9150 29757 9203 29803
rect 9249 29757 9524 29803
rect 9570 29757 9623 29803
rect 9150 29649 9623 29757
rect 9769 29803 10242 29858
rect 9769 29757 9822 29803
rect 9868 29757 10143 29803
rect 10189 29757 10242 29803
rect 9769 29649 10242 29757
rect 10388 29803 10861 29858
rect 10388 29757 10441 29803
rect 10487 29757 10762 29803
rect 10808 29757 10861 29803
rect 10388 29649 10861 29757
rect 11007 29803 11480 29858
rect 11007 29757 11060 29803
rect 11106 29757 11381 29803
rect 11427 29757 11480 29803
rect 11007 29649 11480 29757
rect 11626 29803 12099 29858
rect 11626 29757 11679 29803
rect 11725 29757 12000 29803
rect 12046 29757 12099 29803
rect 11626 29649 12099 29757
rect 12245 29803 12718 29858
rect 12245 29757 12298 29803
rect 12344 29757 12619 29803
rect 12665 29757 12718 29803
rect 12245 29649 12718 29757
rect 12864 29803 13337 29858
rect 12864 29757 12917 29803
rect 12963 29757 13238 29803
rect 13284 29757 13337 29803
rect 12864 29649 13337 29757
rect 13483 29803 13956 29858
rect 13483 29757 13536 29803
rect 13582 29757 13857 29803
rect 13903 29757 13956 29803
rect 13483 29649 13956 29757
rect 14102 29803 14575 29858
rect 14102 29757 14155 29803
rect 14201 29757 14476 29803
rect 14522 29757 14575 29803
rect 14102 29649 14575 29757
rect 14721 29803 15194 29858
rect 14721 29757 14774 29803
rect 14820 29757 15095 29803
rect 15141 29757 15194 29803
rect 14721 29649 15194 29757
rect 15340 29803 15813 29858
rect 15340 29757 15393 29803
rect 15439 29757 15714 29803
rect 15760 29757 15813 29803
rect 15340 29649 15813 29757
rect 15959 29803 16432 29858
rect 15959 29757 16012 29803
rect 16058 29757 16333 29803
rect 16379 29757 16432 29803
rect 15959 29649 16432 29757
rect 16578 29803 17051 29858
rect 16578 29757 16631 29803
rect 16677 29757 16952 29803
rect 16998 29757 17051 29803
rect 16578 29649 17051 29757
rect 17197 29803 17670 29858
rect 17197 29757 17250 29803
rect 17296 29757 17571 29803
rect 17617 29757 17670 29803
rect 17197 29649 17670 29757
rect 17816 29803 18289 29858
rect 17816 29757 17869 29803
rect 17915 29757 18190 29803
rect 18236 29757 18289 29803
rect 17816 29649 18289 29757
rect 18435 29803 18908 29858
rect 18435 29757 18488 29803
rect 18534 29757 18809 29803
rect 18855 29757 18908 29803
rect 18435 29649 18908 29757
rect 19054 29803 19527 29858
rect 19054 29757 19107 29803
rect 19153 29757 19428 29803
rect 19474 29757 19527 29803
rect 19054 29649 19527 29757
rect 19673 29803 20146 29858
rect 19673 29757 19726 29803
rect 19772 29757 20047 29803
rect 20093 29757 20146 29803
rect 19673 29649 20146 29757
rect 20292 29803 20765 29858
rect 20292 29757 20345 29803
rect 20391 29757 20666 29803
rect 20712 29757 20765 29803
rect 20292 29649 20765 29757
rect 20911 29803 21384 29858
rect 20911 29757 20964 29803
rect 21010 29757 21285 29803
rect 21331 29757 21384 29803
rect 20911 29649 21384 29757
rect -754 29112 -281 29194
rect -135 29112 338 29194
rect 484 29112 957 29194
rect 1103 29112 1576 29194
rect 1722 29112 2195 29194
rect 2341 29112 2814 29194
rect 2960 29112 3433 29194
rect 3579 29112 4052 29194
rect 4198 29112 4671 29194
rect 4817 29112 5290 29194
rect 5436 29112 5909 29194
rect 6055 29112 6528 29194
rect 6674 29112 7147 29194
rect 7293 29112 7766 29194
rect 7912 29112 8385 29194
rect 8531 29112 9004 29194
rect 9150 29112 9623 29194
rect 9769 29112 10242 29194
rect 10388 29112 10861 29194
rect 11007 29112 11480 29194
rect 11626 29112 12099 29194
rect 12245 29112 12718 29194
rect 12864 29112 13337 29194
rect 13483 29112 13956 29194
rect 14102 29112 14575 29194
rect 14721 29112 15194 29194
rect 15340 29112 15813 29194
rect 15959 29112 16432 29194
rect 16578 29112 17051 29194
rect 17197 29112 17670 29194
rect 17816 29112 18289 29194
rect 18435 29112 18908 29194
rect 19054 29112 19527 29194
rect 19673 29112 20146 29194
rect 20292 29112 20765 29194
rect 20911 29112 21384 29194
<< polycontact >>
rect -701 29757 -655 29803
rect -380 29757 -334 29803
rect -82 29757 -36 29803
rect 239 29757 285 29803
rect 537 29757 583 29803
rect 858 29757 904 29803
rect 1156 29757 1202 29803
rect 1477 29757 1523 29803
rect 1775 29757 1821 29803
rect 2096 29757 2142 29803
rect 2394 29757 2440 29803
rect 2715 29757 2761 29803
rect 3013 29757 3059 29803
rect 3334 29757 3380 29803
rect 3632 29757 3678 29803
rect 3953 29757 3999 29803
rect 4251 29757 4297 29803
rect 4572 29757 4618 29803
rect 4870 29757 4916 29803
rect 5191 29757 5237 29803
rect 5489 29757 5535 29803
rect 5810 29757 5856 29803
rect 6108 29757 6154 29803
rect 6429 29757 6475 29803
rect 6727 29757 6773 29803
rect 7048 29757 7094 29803
rect 7346 29757 7392 29803
rect 7667 29757 7713 29803
rect 7965 29757 8011 29803
rect 8286 29757 8332 29803
rect 8584 29757 8630 29803
rect 8905 29757 8951 29803
rect 9203 29757 9249 29803
rect 9524 29757 9570 29803
rect 9822 29757 9868 29803
rect 10143 29757 10189 29803
rect 10441 29757 10487 29803
rect 10762 29757 10808 29803
rect 11060 29757 11106 29803
rect 11381 29757 11427 29803
rect 11679 29757 11725 29803
rect 12000 29757 12046 29803
rect 12298 29757 12344 29803
rect 12619 29757 12665 29803
rect 12917 29757 12963 29803
rect 13238 29757 13284 29803
rect 13536 29757 13582 29803
rect 13857 29757 13903 29803
rect 14155 29757 14201 29803
rect 14476 29757 14522 29803
rect 14774 29757 14820 29803
rect 15095 29757 15141 29803
rect 15393 29757 15439 29803
rect 15714 29757 15760 29803
rect 16012 29757 16058 29803
rect 16333 29757 16379 29803
rect 16631 29757 16677 29803
rect 16952 29757 16998 29803
rect 17250 29757 17296 29803
rect 17571 29757 17617 29803
rect 17869 29757 17915 29803
rect 18190 29757 18236 29803
rect 18488 29757 18534 29803
rect 18809 29757 18855 29803
rect 19107 29757 19153 29803
rect 19428 29757 19474 29803
rect 19726 29757 19772 29803
rect 20047 29757 20093 29803
rect 20345 29757 20391 29803
rect 20666 29757 20712 29803
rect 20964 29757 21010 29803
rect 21285 29757 21331 29803
<< metal1 >>
rect -844 29890 -714 30180
rect -1079 29803 21458 29890
rect -1079 29757 -701 29803
rect -655 29757 -380 29803
rect -334 29757 -82 29803
rect -36 29757 239 29803
rect 285 29757 537 29803
rect 583 29757 858 29803
rect 904 29757 1156 29803
rect 1202 29757 1477 29803
rect 1523 29757 1775 29803
rect 1821 29757 2096 29803
rect 2142 29757 2394 29803
rect 2440 29757 2715 29803
rect 2761 29757 3013 29803
rect 3059 29757 3334 29803
rect 3380 29757 3632 29803
rect 3678 29757 3953 29803
rect 3999 29757 4251 29803
rect 4297 29757 4572 29803
rect 4618 29757 4870 29803
rect 4916 29757 5191 29803
rect 5237 29757 5489 29803
rect 5535 29757 5810 29803
rect 5856 29757 6108 29803
rect 6154 29757 6429 29803
rect 6475 29757 6727 29803
rect 6773 29757 7048 29803
rect 7094 29757 7346 29803
rect 7392 29757 7667 29803
rect 7713 29757 7965 29803
rect 8011 29757 8286 29803
rect 8332 29757 8584 29803
rect 8630 29757 8905 29803
rect 8951 29757 9203 29803
rect 9249 29757 9524 29803
rect 9570 29757 9822 29803
rect 9868 29757 10143 29803
rect 10189 29757 10441 29803
rect 10487 29757 10762 29803
rect 10808 29757 11060 29803
rect 11106 29757 11381 29803
rect 11427 29757 11679 29803
rect 11725 29757 12000 29803
rect 12046 29757 12298 29803
rect 12344 29757 12619 29803
rect 12665 29757 12917 29803
rect 12963 29757 13238 29803
rect 13284 29757 13536 29803
rect 13582 29757 13857 29803
rect 13903 29757 14155 29803
rect 14201 29757 14476 29803
rect 14522 29757 14774 29803
rect 14820 29757 15095 29803
rect 15141 29757 15393 29803
rect 15439 29757 15714 29803
rect 15760 29757 16012 29803
rect 16058 29757 16333 29803
rect 16379 29757 16631 29803
rect 16677 29757 16952 29803
rect 16998 29757 17250 29803
rect 17296 29757 17571 29803
rect 17617 29757 17869 29803
rect 17915 29757 18190 29803
rect 18236 29757 18488 29803
rect 18534 29757 18809 29803
rect 18855 29757 19107 29803
rect 19153 29757 19428 29803
rect 19474 29757 19726 29803
rect 19772 29757 20047 29803
rect 20093 29757 20345 29803
rect 20391 29757 20666 29803
rect 20712 29757 20964 29803
rect 21010 29757 21285 29803
rect 21331 29757 21458 29803
rect -1079 29720 21458 29757
rect -885 29604 -769 29640
rect -885 29558 -850 29604
rect -804 29558 -769 29604
rect -885 29286 -769 29558
rect -885 29240 -850 29286
rect -804 29240 -769 29286
rect -885 28890 -769 29240
rect -266 29604 -150 29640
rect -266 29558 -231 29604
rect -185 29558 -150 29604
rect -266 29286 -150 29558
rect -266 29240 -231 29286
rect -185 29240 -150 29286
rect -266 28890 -150 29240
rect 353 29604 469 29640
rect 353 29558 388 29604
rect 434 29558 469 29604
rect 353 29286 469 29558
rect 353 29240 388 29286
rect 434 29240 469 29286
rect 353 28890 469 29240
rect 972 29604 1088 29640
rect 972 29558 1007 29604
rect 1053 29558 1088 29604
rect 972 29286 1088 29558
rect 972 29240 1007 29286
rect 1053 29240 1088 29286
rect 972 28890 1088 29240
rect 1591 29604 1707 29640
rect 1591 29558 1626 29604
rect 1672 29558 1707 29604
rect 1591 29286 1707 29558
rect 1591 29240 1626 29286
rect 1672 29240 1707 29286
rect 1591 28890 1707 29240
rect 2210 29604 2326 29640
rect 2210 29558 2245 29604
rect 2291 29558 2326 29604
rect 2210 29286 2326 29558
rect 2210 29240 2245 29286
rect 2291 29240 2326 29286
rect 2210 28890 2326 29240
rect 2829 29604 2945 29640
rect 2829 29558 2864 29604
rect 2910 29558 2945 29604
rect 2829 29286 2945 29558
rect 2829 29240 2864 29286
rect 2910 29240 2945 29286
rect 2829 28890 2945 29240
rect 3448 29604 3564 29640
rect 3448 29558 3483 29604
rect 3529 29558 3564 29604
rect 3448 29286 3564 29558
rect 3448 29240 3483 29286
rect 3529 29240 3564 29286
rect 3448 28890 3564 29240
rect 4067 29604 4183 29640
rect 4067 29558 4102 29604
rect 4148 29558 4183 29604
rect 4067 29286 4183 29558
rect 4067 29240 4102 29286
rect 4148 29240 4183 29286
rect 4067 28890 4183 29240
rect 4686 29604 4802 29640
rect 4686 29558 4721 29604
rect 4767 29558 4802 29604
rect 4686 29286 4802 29558
rect 4686 29240 4721 29286
rect 4767 29240 4802 29286
rect 4686 28890 4802 29240
rect 5305 29604 5421 29640
rect 5305 29558 5340 29604
rect 5386 29558 5421 29604
rect 5305 29286 5421 29558
rect 5305 29240 5340 29286
rect 5386 29240 5421 29286
rect 5305 28890 5421 29240
rect 5924 29604 6040 29640
rect 5924 29558 5959 29604
rect 6005 29558 6040 29604
rect 5924 29286 6040 29558
rect 5924 29240 5959 29286
rect 6005 29240 6040 29286
rect 5924 28890 6040 29240
rect 6543 29604 6659 29640
rect 6543 29558 6578 29604
rect 6624 29558 6659 29604
rect 6543 29286 6659 29558
rect 6543 29240 6578 29286
rect 6624 29240 6659 29286
rect 6543 28890 6659 29240
rect 7162 29604 7278 29640
rect 7162 29558 7197 29604
rect 7243 29558 7278 29604
rect 7162 29286 7278 29558
rect 7162 29240 7197 29286
rect 7243 29240 7278 29286
rect 7162 28890 7278 29240
rect 7781 29604 7897 29640
rect 7781 29558 7816 29604
rect 7862 29558 7897 29604
rect 7781 29286 7897 29558
rect 7781 29240 7816 29286
rect 7862 29240 7897 29286
rect 7781 28890 7897 29240
rect 8400 29604 8516 29640
rect 8400 29558 8435 29604
rect 8481 29558 8516 29604
rect 8400 29286 8516 29558
rect 8400 29240 8435 29286
rect 8481 29240 8516 29286
rect 8400 28890 8516 29240
rect 9019 29604 9135 29640
rect 9019 29558 9054 29604
rect 9100 29558 9135 29604
rect 9019 29286 9135 29558
rect 9019 29240 9054 29286
rect 9100 29240 9135 29286
rect 9019 28890 9135 29240
rect 9638 29604 9754 29640
rect 9638 29558 9673 29604
rect 9719 29558 9754 29604
rect 9638 29286 9754 29558
rect 9638 29240 9673 29286
rect 9719 29240 9754 29286
rect 9638 28890 9754 29240
rect 10257 29604 10373 29640
rect 10257 29558 10292 29604
rect 10338 29558 10373 29604
rect 10257 29286 10373 29558
rect 10257 29240 10292 29286
rect 10338 29240 10373 29286
rect 10257 28890 10373 29240
rect 10876 29604 10992 29640
rect 10876 29558 10911 29604
rect 10957 29558 10992 29604
rect 10876 29286 10992 29558
rect 10876 29240 10911 29286
rect 10957 29240 10992 29286
rect 10876 28890 10992 29240
rect 11495 29604 11611 29640
rect 11495 29558 11530 29604
rect 11576 29558 11611 29604
rect 11495 29286 11611 29558
rect 11495 29240 11530 29286
rect 11576 29240 11611 29286
rect 11495 28890 11611 29240
rect 12114 29604 12230 29640
rect 12114 29558 12149 29604
rect 12195 29558 12230 29604
rect 12114 29286 12230 29558
rect 12114 29240 12149 29286
rect 12195 29240 12230 29286
rect 12114 28890 12230 29240
rect 12733 29604 12849 29640
rect 12733 29558 12768 29604
rect 12814 29558 12849 29604
rect 12733 29286 12849 29558
rect 12733 29240 12768 29286
rect 12814 29240 12849 29286
rect 12733 28890 12849 29240
rect 13352 29604 13468 29640
rect 13352 29558 13387 29604
rect 13433 29558 13468 29604
rect 13352 29286 13468 29558
rect 13352 29240 13387 29286
rect 13433 29240 13468 29286
rect 13352 28890 13468 29240
rect 13971 29604 14087 29640
rect 13971 29558 14006 29604
rect 14052 29558 14087 29604
rect 13971 29286 14087 29558
rect 13971 29240 14006 29286
rect 14052 29240 14087 29286
rect 13971 28890 14087 29240
rect 14590 29604 14706 29640
rect 14590 29558 14625 29604
rect 14671 29558 14706 29604
rect 14590 29286 14706 29558
rect 14590 29240 14625 29286
rect 14671 29240 14706 29286
rect 14590 28890 14706 29240
rect 15209 29604 15325 29640
rect 15209 29558 15244 29604
rect 15290 29558 15325 29604
rect 15209 29286 15325 29558
rect 15209 29240 15244 29286
rect 15290 29240 15325 29286
rect 15209 28890 15325 29240
rect 15828 29604 15944 29640
rect 15828 29558 15863 29604
rect 15909 29558 15944 29604
rect 15828 29286 15944 29558
rect 15828 29240 15863 29286
rect 15909 29240 15944 29286
rect 15828 28890 15944 29240
rect 16447 29604 16563 29640
rect 16447 29558 16482 29604
rect 16528 29558 16563 29604
rect 16447 29286 16563 29558
rect 16447 29240 16482 29286
rect 16528 29240 16563 29286
rect 16447 28890 16563 29240
rect 17066 29604 17182 29640
rect 17066 29558 17101 29604
rect 17147 29558 17182 29604
rect 17066 29286 17182 29558
rect 17066 29240 17101 29286
rect 17147 29240 17182 29286
rect 17066 28890 17182 29240
rect 17685 29604 17801 29640
rect 17685 29558 17720 29604
rect 17766 29558 17801 29604
rect 17685 29286 17801 29558
rect 17685 29240 17720 29286
rect 17766 29240 17801 29286
rect 17685 28890 17801 29240
rect 18304 29604 18420 29640
rect 18304 29558 18339 29604
rect 18385 29558 18420 29604
rect 18304 29286 18420 29558
rect 18304 29240 18339 29286
rect 18385 29240 18420 29286
rect 18304 28890 18420 29240
rect 18923 29604 19039 29640
rect 18923 29558 18958 29604
rect 19004 29558 19039 29604
rect 18923 29286 19039 29558
rect 18923 29240 18958 29286
rect 19004 29240 19039 29286
rect 18923 28890 19039 29240
rect 19542 29604 19658 29640
rect 19542 29558 19577 29604
rect 19623 29558 19658 29604
rect 19542 29286 19658 29558
rect 19542 29240 19577 29286
rect 19623 29240 19658 29286
rect 19542 28890 19658 29240
rect 20161 29604 20277 29640
rect 20161 29558 20196 29604
rect 20242 29558 20277 29604
rect 20161 29286 20277 29558
rect 20161 29240 20196 29286
rect 20242 29240 20277 29286
rect 20161 28890 20277 29240
rect 20780 29604 20896 29640
rect 20780 29558 20815 29604
rect 20861 29558 20896 29604
rect 20780 29286 20896 29558
rect 20780 29240 20815 29286
rect 20861 29240 20896 29286
rect 20780 28890 20896 29240
rect 21399 29604 21515 29640
rect 21399 29558 21434 29604
rect 21480 29558 21515 29604
rect 21399 29286 21515 29558
rect 21399 29240 21434 29286
rect 21480 29240 21515 29286
rect 21399 28890 21515 29240
rect -885 28725 21515 28890
<< metal2 >>
rect -827 29107 -738 29955
rect -827 29069 -733 29107
rect -827 29013 -808 29069
rect -752 29013 -733 29069
rect -827 28883 -733 29013
rect -827 28827 -808 28883
rect -752 28827 -733 28883
rect -827 28788 -733 28827
rect -827 21746 -738 28788
<< via2 >>
rect -808 29013 -752 29069
rect -808 28827 -752 28883
<< metal3 >>
rect -1115 88917 21718 89277
rect -1059 40473 -831 40623
rect -1 29713 640 29846
rect -826 29069 -733 29107
rect -826 29013 -808 29069
rect -752 29013 -733 29069
rect -826 28883 -733 29013
rect -826 28827 -808 28883
rect -752 28827 -733 28883
rect -826 28788 -733 28827
use col_512a_512x8m81  col_512a_512x8m81_0
timestamp 1750858719
transform 1 0 -13 0 1 -1433
box -1222 -1965 22823 90208
use dcap_103_novia_512x8m81  dcap_103_novia_512x8m81_0
array 0 35 619 0 0 0
timestamp 1750858719
transform 1 0 -827 0 1 29009
box 0 0 1 1
use ldummy_512x4_512x8m81  ldummy_512x4_512x8m81_0
timestamp 1750858719
transform 1 0 -541 0 1 30030
box -636 76 22573 59677
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1750858719
transform 1 0 -826 0 1 28789
box 0 0 1 1
<< labels >>
rlabel metal3 s 685 60366 685 60366 4 WL[32]
port 1 nsew
rlabel metal3 s 685 61266 685 61266 4 WL[33]
port 2 nsew
rlabel metal3 s 685 62166 685 62166 4 WL[34]
port 3 nsew
rlabel metal3 s 685 65766 685 65766 4 WL[38]
port 4 nsew
rlabel metal3 s 685 66666 685 66666 4 WL[39]
port 5 nsew
rlabel metal3 s 685 63066 685 63066 4 WL[35]
port 6 nsew
rlabel metal3 s 685 63966 685 63966 4 WL[36]
port 7 nsew
rlabel metal3 s 685 64866 685 64866 4 WL[37]
port 8 nsew
rlabel metal3 s 685 67566 685 67566 4 WL[40]
port 9 nsew
rlabel metal3 s 685 68466 685 68466 4 WL[41]
port 10 nsew
rlabel metal3 s 685 69366 685 69366 4 WL[42]
port 11 nsew
rlabel metal3 s 685 70266 685 70266 4 WL[43]
port 12 nsew
rlabel metal3 s 685 71166 685 71166 4 WL[44]
port 13 nsew
rlabel metal3 s 685 72066 685 72066 4 WL[45]
port 14 nsew
rlabel metal3 s 685 72966 685 72966 4 WL[46]
port 15 nsew
rlabel metal3 s 685 73866 685 73866 4 WL[47]
port 16 nsew
rlabel metal3 s 685 74766 685 74766 4 WL[48]
port 17 nsew
rlabel metal3 s 685 75666 685 75666 4 WL[49]
port 18 nsew
rlabel metal3 s 685 76566 685 76566 4 WL[50]
port 19 nsew
rlabel metal3 s 685 77466 685 77466 4 WL[51]
port 20 nsew
rlabel metal3 s 685 78366 685 78366 4 WL[52]
port 21 nsew
rlabel metal3 s 685 79266 685 79266 4 WL[53]
port 22 nsew
rlabel metal3 s 685 80166 685 80166 4 WL[54]
port 23 nsew
rlabel metal3 s 685 81066 685 81066 4 WL[55]
port 24 nsew
rlabel metal3 s 685 81966 685 81966 4 WL[56]
port 25 nsew
rlabel metal3 s 685 82866 685 82866 4 WL[57]
port 26 nsew
rlabel metal3 s 685 83766 685 83766 4 WL[58]
port 27 nsew
rlabel metal3 s 685 84666 685 84666 4 WL[59]
port 28 nsew
rlabel metal3 s 685 85566 685 85566 4 WL[60]
port 29 nsew
rlabel metal3 s 685 86466 685 86466 4 WL[61]
port 30 nsew
rlabel metal3 s 685 87366 685 87366 4 WL[62]
port 31 nsew
rlabel metal3 s 685 88266 685 88266 4 WL[63]
port 32 nsew
rlabel metal3 s 701 54068 701 54068 4 WL[25]
port 33 nsew
rlabel metal3 s 701 53168 701 53168 4 WL[24]
port 34 nsew
rlabel metal3 s 701 52268 701 52268 4 WL[23]
port 35 nsew
rlabel metal3 s 701 51368 701 51368 4 WL[22]
port 36 nsew
rlabel metal3 s 701 50468 701 50468 4 WL[21]
port 37 nsew
rlabel metal3 s 701 49568 701 49568 4 WL[20]
port 38 nsew
rlabel metal3 s 701 48668 701 48668 4 WL[19]
port 39 nsew
rlabel metal3 s 701 47768 701 47768 4 WL[18]
port 40 nsew
rlabel metal3 s 701 46868 701 46868 4 WL[17]
port 41 nsew
rlabel metal3 s 701 45968 701 45968 4 WL[16]
port 42 nsew
rlabel metal3 s 701 45068 701 45068 4 WL[15]
port 43 nsew
rlabel metal3 s 701 44168 701 44168 4 WL[14]
port 44 nsew
rlabel metal3 s 701 43268 701 43268 4 WL[13]
port 45 nsew
rlabel metal3 s 701 42368 701 42368 4 WL[12]
port 46 nsew
rlabel metal3 s 701 41468 701 41468 4 WL[11]
port 47 nsew
rlabel metal3 s 701 40568 701 40568 4 WL[10]
port 48 nsew
rlabel metal3 s 701 39668 701 39668 4 WL[9]
port 49 nsew
rlabel metal3 s 701 38768 701 38768 4 WL[8]
port 50 nsew
rlabel metal3 s 701 37868 701 37868 4 WL[7]
port 51 nsew
rlabel metal3 s 701 36968 701 36968 4 WL[6]
port 52 nsew
rlabel metal3 s 701 36068 701 36068 4 WL[5]
port 53 nsew
rlabel metal3 s 701 35168 701 35168 4 WL[4]
port 54 nsew
rlabel metal3 s 701 34268 701 34268 4 WL[3]
port 55 nsew
rlabel metal3 s 701 33368 701 33368 4 WL[2]
port 56 nsew
rlabel metal3 s 701 32468 701 32468 4 WL[1]
port 57 nsew
rlabel metal3 s 701 31568 701 31568 4 WL[0]
port 58 nsew
rlabel metal3 s 701 59468 701 59468 4 WL[31]
port 59 nsew
rlabel metal3 s 701 58568 701 58568 4 WL[30]
port 60 nsew
rlabel metal3 s 701 57668 701 57668 4 WL[29]
port 61 nsew
rlabel metal3 s 701 56768 701 56768 4 WL[28]
port 62 nsew
rlabel metal3 s 701 55868 701 55868 4 WL[27]
port 63 nsew
rlabel metal3 s 701 54968 701 54968 4 WL[26]
port 64 nsew
rlabel metal3 s 870 1467 870 1467 4 men
port 65 nsew
rlabel metal3 s 797 18592 797 18592 4 ypass[0]
port 66 nsew
rlabel metal3 s 797 18914 797 18914 4 ypass[1]
port 67 nsew
rlabel metal3 s 797 19231 797 19231 4 ypass[2]
port 68 nsew
rlabel metal3 s 797 19548 797 19548 4 ypass[3]
port 69 nsew
rlabel metal3 s 797 20204 797 20204 4 ypass[4]
port 70 nsew
rlabel metal3 s 797 20528 797 20528 4 ypass[5]
port 71 nsew
rlabel metal3 s 797 20845 797 20845 4 ypass[6]
port 72 nsew
rlabel metal3 s 797 21162 797 21162 4 ypass[7]
port 73 nsew
rlabel metal3 s 867 1467 867 1467 4 men
port 65 nsew
flabel metal3 s -334 8814 -334 8814 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 386 -334 386 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -305 1002 -305 1002 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 2322 -305 2322 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 5923 -305 5923 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 11468 -305 11468 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 17107 -305 17107 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 22970 -305 22970 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 29782 -305 29782 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -334 3858 -334 3858 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 7580 -334 7580 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 14009 -334 14009 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 18141 -334 18141 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 27925 -334 27925 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 -708 -334 -708 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -334 -3027 -334 -3027 0 FreeSans 1600 0 0 0 VDD
port 74 nsew
flabel metal3 s -305 -1478 -305 -1478 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s -305 -2341 -305 -2341 0 FreeSans 1600 0 0 0 VSS
port 75 nsew
flabel metal3 s 793 -1999 793 -1999 0 FreeSans 1600 0 0 0 GWEN
port 76 nsew
flabel metal3 s -325 4973 -325 4973 0 FreeSans 1600 0 0 0 GWE
port 77 nsew
rlabel metal2 s -477 104 -477 104 4 din[0]
port 78 nsew
rlabel metal2 s 9695 104 9695 104 4 din[1]
port 79 nsew
rlabel metal2 s 20487 104 20487 104 4 din[3]
port 80 nsew
rlabel metal2 s 10332 104 10332 104 4 din[2]
port 81 nsew
rlabel metal2 s 370 104 370 104 4 q[0]
port 82 nsew
rlabel metal2 s 8853 104 8853 104 4 q[1]
port 83 nsew
rlabel metal2 s 11190 104 11190 104 4 q[2]
port 84 nsew
rlabel metal2 s 19651 104 19651 104 4 q[3]
port 85 nsew
rlabel metal1 s 5690 15928 5690 15928 4 pcb[2]
port 86 nsew
rlabel metal1 s 3660 15928 3660 15928 4 pcb[3]
port 87 nsew
rlabel metal1 s 16496 15928 16496 15928 4 pcb[0]
port 88 nsew
rlabel metal1 s 14155 15928 14155 15928 4 pcb[1]
port 89 nsew
rlabel metal1 s 920 18163 920 18163 4 vdd
port 90 nsew
flabel metal1 s -808 31106 -808 31106 0 FreeSans 368 0 0 0 VDD
port 74 nsew
flabel metal1 s -367 -3355 -367 -3355 0 FreeSans 600 0 0 0 WEN[3]
port 91 nsew
flabel metal1 s 9597 -3329 9597 -3329 0 FreeSans 600 0 0 0 WEN[2]
port 92 nsew
flabel metal1 s 10395 -3329 10395 -3329 0 FreeSans 600 0 0 0 WEN[1]
port 93 nsew
flabel metal1 s 20398 -3329 20398 -3329 0 FreeSans 600 0 0 0 WEN[0]
port 94 nsew
<< properties >>
string GDS_END 2648100
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2641714
<< end >>
