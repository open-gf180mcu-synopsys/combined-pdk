magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< isosubstrate >>
rect 2248 55601 14818 56937
rect 4664 55565 7604 55601
rect 9908 55565 12848 55601
rect 10564 42246 14743 43312
rect 11970 40612 14743 42246
<< nwell >>
rect 955 54474 2177 55927
rect 873 52942 2754 54474
rect 11242 40577 11874 41673
<< pwell >>
rect 2760 56031 3760 56507
rect 4260 56031 5260 56507
rect 5760 56031 6760 56507
rect 7260 56031 8260 56507
rect 8760 56031 9760 56507
rect 10260 56031 11260 56507
rect 11760 56031 12760 56507
rect 13260 56031 14260 56507
rect 12482 42058 13082 42834
rect 13622 42058 14222 42834
rect 12482 41090 13082 41866
rect 13622 41090 14222 41866
<< mvndiff >>
rect 2760 56494 3760 56507
rect 2760 56448 2797 56494
rect 3723 56448 3760 56494
rect 2760 56419 3760 56448
rect 4260 56494 5260 56507
rect 4260 56448 4297 56494
rect 5223 56448 5260 56494
rect 4260 56419 5260 56448
rect 5760 56494 6760 56507
rect 5760 56448 5797 56494
rect 6723 56448 6760 56494
rect 5760 56419 6760 56448
rect 7260 56494 8260 56507
rect 7260 56448 7297 56494
rect 8223 56448 8260 56494
rect 7260 56419 8260 56448
rect 8760 56494 9760 56507
rect 8760 56448 8797 56494
rect 9723 56448 9760 56494
rect 8760 56419 9760 56448
rect 10260 56494 11260 56507
rect 10260 56448 10297 56494
rect 11223 56448 11260 56494
rect 10260 56419 11260 56448
rect 11760 56494 12760 56507
rect 11760 56448 11797 56494
rect 12723 56448 12760 56494
rect 11760 56419 12760 56448
rect 13260 56494 14260 56507
rect 13260 56448 13297 56494
rect 14223 56448 14260 56494
rect 13260 56419 14260 56448
rect 2760 56090 3760 56119
rect 2760 56044 2797 56090
rect 3723 56044 3760 56090
rect 2760 56031 3760 56044
rect 4260 56090 5260 56119
rect 4260 56044 4297 56090
rect 5223 56044 5260 56090
rect 4260 56031 5260 56044
rect 5760 56090 6760 56119
rect 5760 56044 5797 56090
rect 6723 56044 6760 56090
rect 5760 56031 6760 56044
rect 7260 56090 8260 56119
rect 7260 56044 7297 56090
rect 8223 56044 8260 56090
rect 7260 56031 8260 56044
rect 8760 56090 9760 56119
rect 8760 56044 8797 56090
rect 9723 56044 9760 56090
rect 8760 56031 9760 56044
rect 10260 56090 11260 56119
rect 10260 56044 10297 56090
rect 11223 56044 11260 56090
rect 10260 56031 11260 56044
rect 11760 56090 12760 56119
rect 11760 56044 11797 56090
rect 12723 56044 12760 56090
rect 11760 56031 12760 56044
rect 13260 56090 14260 56119
rect 13260 56044 13297 56090
rect 14223 56044 14260 56090
rect 13260 56031 14260 56044
rect 12482 42821 13082 42834
rect 12482 42775 12519 42821
rect 13045 42775 13082 42821
rect 12482 42746 13082 42775
rect 13622 42821 14222 42834
rect 13622 42775 13659 42821
rect 14185 42775 14222 42821
rect 13622 42746 14222 42775
rect 12482 42117 13082 42146
rect 12482 42071 12519 42117
rect 13045 42071 13082 42117
rect 12482 42058 13082 42071
rect 13622 42117 14222 42146
rect 13622 42071 13659 42117
rect 14185 42071 14222 42117
rect 13622 42058 14222 42071
rect 12482 41853 13082 41866
rect 12482 41807 12519 41853
rect 13045 41807 13082 41853
rect 12482 41778 13082 41807
rect 13622 41853 14222 41866
rect 13622 41807 13659 41853
rect 14185 41807 14222 41853
rect 13622 41778 14222 41807
rect 12482 41149 13082 41178
rect 12482 41103 12519 41149
rect 13045 41103 13082 41149
rect 12482 41090 13082 41103
rect 13622 41149 14222 41178
rect 13622 41103 13659 41149
rect 14185 41103 14222 41149
rect 13622 41090 14222 41103
<< mvndiffc >>
rect 2797 56448 3723 56494
rect 4297 56448 5223 56494
rect 5797 56448 6723 56494
rect 7297 56448 8223 56494
rect 8797 56448 9723 56494
rect 10297 56448 11223 56494
rect 11797 56448 12723 56494
rect 13297 56448 14223 56494
rect 2797 56044 3723 56090
rect 4297 56044 5223 56090
rect 5797 56044 6723 56090
rect 7297 56044 8223 56090
rect 8797 56044 9723 56090
rect 10297 56044 11223 56090
rect 11797 56044 12723 56090
rect 13297 56044 14223 56090
rect 12519 42775 13045 42821
rect 13659 42775 14185 42821
rect 12519 42071 13045 42117
rect 13659 42071 14185 42117
rect 12519 41807 13045 41853
rect 13659 41807 14185 41853
rect 12519 41103 13045 41149
rect 13659 41103 14185 41149
<< psubdiff >>
rect 2331 56832 14735 56854
rect 2331 56786 2353 56832
rect 14713 56786 14735 56832
rect 2331 56764 14735 56786
rect 2331 56668 2421 56764
rect 2331 55870 2353 56668
rect 2399 55870 2421 56668
rect 14645 56668 14735 56764
rect 2331 55774 2421 55870
rect 14645 55870 14667 56668
rect 14713 55870 14735 56668
rect 14645 55774 14735 55870
rect 2331 55752 14735 55774
rect 2331 55706 2353 55752
rect 14713 55706 14735 55752
rect 2331 55684 14735 55706
rect 10742 43258 11858 43280
rect 10742 43212 10764 43258
rect 10810 43212 10878 43258
rect 10924 43212 10992 43258
rect 11038 43212 11106 43258
rect 11152 43212 11220 43258
rect 11266 43212 11334 43258
rect 11380 43212 11448 43258
rect 11494 43212 11562 43258
rect 11608 43212 11676 43258
rect 11722 43212 11790 43258
rect 11836 43212 11858 43258
rect 10742 43144 11858 43212
rect 10742 43098 10764 43144
rect 10810 43098 10878 43144
rect 10924 43098 10992 43144
rect 11038 43098 11106 43144
rect 11152 43098 11220 43144
rect 11266 43098 11334 43144
rect 11380 43098 11448 43144
rect 11494 43098 11562 43144
rect 11608 43098 11676 43144
rect 11722 43098 11790 43144
rect 11836 43098 11858 43144
rect 10742 43030 11858 43098
rect 10742 42984 10764 43030
rect 10810 42984 10878 43030
rect 10924 42984 10992 43030
rect 11038 42984 11106 43030
rect 11152 42984 11220 43030
rect 11266 42984 11334 43030
rect 11380 42984 11448 43030
rect 11494 42984 11562 43030
rect 11608 42984 11676 43030
rect 11722 42984 11790 43030
rect 11836 42984 11858 43030
rect 10742 42916 11858 42984
rect 10742 42870 10764 42916
rect 10810 42870 10878 42916
rect 10924 42870 10992 42916
rect 11038 42870 11106 42916
rect 11152 42870 11220 42916
rect 11266 42870 11334 42916
rect 11380 42870 11448 42916
rect 11494 42870 11562 42916
rect 11608 42870 11676 42916
rect 11722 42870 11790 42916
rect 11836 42870 11858 42916
rect 10742 42802 11858 42870
rect 10742 42756 10764 42802
rect 10810 42756 10878 42802
rect 10924 42756 10992 42802
rect 11038 42756 11106 42802
rect 11152 42756 11220 42802
rect 11266 42756 11334 42802
rect 11380 42756 11448 42802
rect 11494 42756 11562 42802
rect 11608 42756 11676 42802
rect 11722 42756 11790 42802
rect 11836 42756 11858 42802
rect 10742 42688 11858 42756
rect 10742 42642 10764 42688
rect 10810 42642 10878 42688
rect 10924 42642 10992 42688
rect 11038 42642 11106 42688
rect 11152 42642 11220 42688
rect 11266 42642 11334 42688
rect 11380 42642 11448 42688
rect 11494 42642 11562 42688
rect 11608 42642 11676 42688
rect 11722 42642 11790 42688
rect 11836 42642 11858 42688
rect 10742 42574 11858 42642
rect 10742 42528 10764 42574
rect 10810 42528 10878 42574
rect 10924 42528 10992 42574
rect 11038 42528 11106 42574
rect 11152 42528 11220 42574
rect 11266 42528 11334 42574
rect 11380 42528 11448 42574
rect 11494 42528 11562 42574
rect 11608 42528 11676 42574
rect 11722 42528 11790 42574
rect 11836 42528 11858 42574
rect 10742 42460 11858 42528
rect 10742 42414 10764 42460
rect 10810 42414 10878 42460
rect 10924 42414 10992 42460
rect 11038 42414 11106 42460
rect 11152 42414 11220 42460
rect 11266 42414 11334 42460
rect 11380 42414 11448 42460
rect 11494 42414 11562 42460
rect 11608 42414 11676 42460
rect 11722 42414 11790 42460
rect 11836 42414 11858 42460
rect 10742 42346 11858 42414
rect 10742 42300 10764 42346
rect 10810 42300 10878 42346
rect 10924 42300 10992 42346
rect 11038 42300 11106 42346
rect 11152 42300 11220 42346
rect 11266 42300 11334 42346
rect 11380 42300 11448 42346
rect 11494 42300 11562 42346
rect 11608 42300 11676 42346
rect 11722 42300 11790 42346
rect 11836 42300 11858 42346
rect 10742 42278 11858 42300
rect 12053 43207 14660 43229
rect 12053 40717 12075 43207
rect 12121 43161 12182 43207
rect 14484 43161 14592 43207
rect 12121 43139 14592 43161
rect 12121 40785 12143 43139
rect 14570 40785 14592 43139
rect 12121 40763 14592 40785
rect 12121 40717 12182 40763
rect 14484 40717 14592 40763
rect 14638 40717 14660 43207
rect 12053 40695 14660 40717
rect 257 9265 843 9287
rect 257 9219 279 9265
rect 325 9219 403 9265
rect 449 9219 527 9265
rect 573 9219 651 9265
rect 697 9219 775 9265
rect 821 9219 843 9265
rect 257 9141 843 9219
rect 257 9095 279 9141
rect 325 9095 403 9141
rect 449 9095 527 9141
rect 573 9095 651 9141
rect 697 9095 775 9141
rect 821 9095 843 9141
rect 257 9017 843 9095
rect 257 8971 279 9017
rect 325 8971 403 9017
rect 449 8971 527 9017
rect 573 8971 651 9017
rect 697 8971 775 9017
rect 821 8971 843 9017
rect 257 8893 843 8971
rect 257 8847 279 8893
rect 325 8847 403 8893
rect 449 8847 527 8893
rect 573 8847 651 8893
rect 697 8847 775 8893
rect 821 8847 843 8893
rect 257 8769 843 8847
rect 257 8723 279 8769
rect 325 8723 403 8769
rect 449 8723 527 8769
rect 573 8723 651 8769
rect 697 8723 775 8769
rect 821 8723 843 8769
rect 257 8645 843 8723
rect 257 8599 279 8645
rect 325 8599 403 8645
rect 449 8599 527 8645
rect 573 8599 651 8645
rect 697 8599 775 8645
rect 821 8599 843 8645
rect 257 8521 843 8599
rect 257 8475 279 8521
rect 325 8475 403 8521
rect 449 8475 527 8521
rect 573 8475 651 8521
rect 697 8475 775 8521
rect 821 8475 843 8521
rect 257 8397 843 8475
rect 257 8351 279 8397
rect 325 8351 403 8397
rect 449 8351 527 8397
rect 573 8351 651 8397
rect 697 8351 775 8397
rect 821 8351 843 8397
rect 257 8273 843 8351
rect 257 8227 279 8273
rect 325 8227 403 8273
rect 449 8227 527 8273
rect 573 8227 651 8273
rect 697 8227 775 8273
rect 821 8227 843 8273
rect 257 8149 843 8227
rect 257 8103 279 8149
rect 325 8103 403 8149
rect 449 8103 527 8149
rect 573 8103 651 8149
rect 697 8103 775 8149
rect 821 8103 843 8149
rect 257 8025 843 8103
rect 257 7979 279 8025
rect 325 7979 403 8025
rect 449 7979 527 8025
rect 573 7979 651 8025
rect 697 7979 775 8025
rect 821 7979 843 8025
rect 257 7901 843 7979
rect 257 7855 279 7901
rect 325 7855 403 7901
rect 449 7855 527 7901
rect 573 7855 651 7901
rect 697 7855 775 7901
rect 821 7855 843 7901
rect 257 7777 843 7855
rect 257 7731 279 7777
rect 325 7731 403 7777
rect 449 7731 527 7777
rect 573 7731 651 7777
rect 697 7731 775 7777
rect 821 7731 843 7777
rect 257 7653 843 7731
rect 257 7607 279 7653
rect 325 7607 403 7653
rect 449 7607 527 7653
rect 573 7607 651 7653
rect 697 7607 775 7653
rect 821 7607 843 7653
rect 257 7529 843 7607
rect 257 7483 279 7529
rect 325 7483 403 7529
rect 449 7483 527 7529
rect 573 7483 651 7529
rect 697 7483 775 7529
rect 821 7483 843 7529
rect 257 7405 843 7483
rect 257 7359 279 7405
rect 325 7359 403 7405
rect 449 7359 527 7405
rect 573 7359 651 7405
rect 697 7359 775 7405
rect 821 7359 843 7405
rect 257 7281 843 7359
rect 257 7235 279 7281
rect 325 7235 403 7281
rect 449 7235 527 7281
rect 573 7235 651 7281
rect 697 7235 775 7281
rect 821 7235 843 7281
rect 257 7157 843 7235
rect 257 7111 279 7157
rect 325 7111 403 7157
rect 449 7111 527 7157
rect 573 7111 651 7157
rect 697 7111 775 7157
rect 821 7111 843 7157
rect 257 7033 843 7111
rect 257 6987 279 7033
rect 325 6987 403 7033
rect 449 6987 527 7033
rect 573 6987 651 7033
rect 697 6987 775 7033
rect 821 6987 843 7033
rect 257 6909 843 6987
rect 257 6863 279 6909
rect 325 6863 403 6909
rect 449 6863 527 6909
rect 573 6863 651 6909
rect 697 6863 775 6909
rect 821 6863 843 6909
rect 257 6785 843 6863
rect 257 6739 279 6785
rect 325 6739 403 6785
rect 449 6739 527 6785
rect 573 6739 651 6785
rect 697 6739 775 6785
rect 821 6739 843 6785
rect 257 6661 843 6739
rect 257 6615 279 6661
rect 325 6615 403 6661
rect 449 6615 527 6661
rect 573 6615 651 6661
rect 697 6615 775 6661
rect 821 6615 843 6661
rect 257 6537 843 6615
rect 257 6491 279 6537
rect 325 6491 403 6537
rect 449 6491 527 6537
rect 573 6491 651 6537
rect 697 6491 775 6537
rect 821 6491 843 6537
rect 257 6413 843 6491
rect 257 6367 279 6413
rect 325 6367 403 6413
rect 449 6367 527 6413
rect 573 6367 651 6413
rect 697 6367 775 6413
rect 821 6367 843 6413
rect 257 6289 843 6367
rect 257 6243 279 6289
rect 325 6243 403 6289
rect 449 6243 527 6289
rect 573 6243 651 6289
rect 697 6243 775 6289
rect 821 6243 843 6289
rect 257 6165 843 6243
rect 257 6119 279 6165
rect 325 6119 403 6165
rect 449 6119 527 6165
rect 573 6119 651 6165
rect 697 6119 775 6165
rect 821 6119 843 6165
rect 257 6041 843 6119
rect 257 5995 279 6041
rect 325 5995 403 6041
rect 449 5995 527 6041
rect 573 5995 651 6041
rect 697 5995 775 6041
rect 821 5995 843 6041
rect 257 5917 843 5995
rect 257 5871 279 5917
rect 325 5871 403 5917
rect 449 5871 527 5917
rect 573 5871 651 5917
rect 697 5871 775 5917
rect 821 5871 843 5917
rect 257 5793 843 5871
rect 257 5747 279 5793
rect 325 5747 403 5793
rect 449 5747 527 5793
rect 573 5747 651 5793
rect 697 5747 775 5793
rect 821 5747 843 5793
rect 257 5669 843 5747
rect 257 5623 279 5669
rect 325 5623 403 5669
rect 449 5623 527 5669
rect 573 5623 651 5669
rect 697 5623 775 5669
rect 821 5623 843 5669
rect 257 5545 843 5623
rect 257 5499 279 5545
rect 325 5499 403 5545
rect 449 5499 527 5545
rect 573 5499 651 5545
rect 697 5499 775 5545
rect 821 5499 843 5545
rect 257 5421 843 5499
rect 257 5375 279 5421
rect 325 5375 403 5421
rect 449 5375 527 5421
rect 573 5375 651 5421
rect 697 5375 775 5421
rect 821 5375 843 5421
rect 257 5297 843 5375
rect 257 5251 279 5297
rect 325 5251 403 5297
rect 449 5251 527 5297
rect 573 5251 651 5297
rect 697 5251 775 5297
rect 821 5251 843 5297
rect 257 5173 843 5251
rect 257 5127 279 5173
rect 325 5127 403 5173
rect 449 5127 527 5173
rect 573 5127 651 5173
rect 697 5127 775 5173
rect 821 5127 843 5173
rect 257 5049 843 5127
rect 257 5003 279 5049
rect 325 5003 403 5049
rect 449 5003 527 5049
rect 573 5003 651 5049
rect 697 5003 775 5049
rect 821 5003 843 5049
rect 257 4925 843 5003
rect 257 4879 279 4925
rect 325 4879 403 4925
rect 449 4879 527 4925
rect 573 4879 651 4925
rect 697 4879 775 4925
rect 821 4879 843 4925
rect 257 4801 843 4879
rect 257 4755 279 4801
rect 325 4755 403 4801
rect 449 4755 527 4801
rect 573 4755 651 4801
rect 697 4755 775 4801
rect 821 4755 843 4801
rect 257 4677 843 4755
rect 257 4631 279 4677
rect 325 4631 403 4677
rect 449 4631 527 4677
rect 573 4631 651 4677
rect 697 4631 775 4677
rect 821 4631 843 4677
rect 257 4553 843 4631
rect 257 4507 279 4553
rect 325 4507 403 4553
rect 449 4507 527 4553
rect 573 4507 651 4553
rect 697 4507 775 4553
rect 821 4507 843 4553
rect 257 4429 843 4507
rect 257 4383 279 4429
rect 325 4383 403 4429
rect 449 4383 527 4429
rect 573 4383 651 4429
rect 697 4383 775 4429
rect 821 4383 843 4429
rect 257 4305 843 4383
rect 257 4259 279 4305
rect 325 4259 403 4305
rect 449 4259 527 4305
rect 573 4259 651 4305
rect 697 4259 775 4305
rect 821 4259 843 4305
rect 257 4181 843 4259
rect 257 4135 279 4181
rect 325 4135 403 4181
rect 449 4135 527 4181
rect 573 4135 651 4181
rect 697 4135 775 4181
rect 821 4135 843 4181
rect 257 4057 843 4135
rect 257 4011 279 4057
rect 325 4011 403 4057
rect 449 4011 527 4057
rect 573 4011 651 4057
rect 697 4011 775 4057
rect 821 4011 843 4057
rect 257 3933 843 4011
rect 257 3887 279 3933
rect 325 3887 403 3933
rect 449 3887 527 3933
rect 573 3887 651 3933
rect 697 3887 775 3933
rect 821 3887 843 3933
rect 257 3809 843 3887
rect 257 3763 279 3809
rect 325 3763 403 3809
rect 449 3763 527 3809
rect 573 3763 651 3809
rect 697 3763 775 3809
rect 821 3763 843 3809
rect 257 3685 843 3763
rect 257 3639 279 3685
rect 325 3639 403 3685
rect 449 3639 527 3685
rect 573 3639 651 3685
rect 697 3639 775 3685
rect 821 3639 843 3685
rect 257 3561 843 3639
rect 257 3515 279 3561
rect 325 3515 403 3561
rect 449 3515 527 3561
rect 573 3515 651 3561
rect 697 3515 775 3561
rect 821 3515 843 3561
rect 257 3437 843 3515
rect 257 3391 279 3437
rect 325 3391 403 3437
rect 449 3391 527 3437
rect 573 3391 651 3437
rect 697 3391 775 3437
rect 821 3391 843 3437
rect 257 3313 843 3391
rect 257 3267 279 3313
rect 325 3267 403 3313
rect 449 3267 527 3313
rect 573 3267 651 3313
rect 697 3267 775 3313
rect 821 3267 843 3313
rect 257 3189 843 3267
rect 257 3143 279 3189
rect 325 3143 403 3189
rect 449 3143 527 3189
rect 573 3143 651 3189
rect 697 3143 775 3189
rect 821 3143 843 3189
rect 257 3065 843 3143
rect 257 3019 279 3065
rect 325 3019 403 3065
rect 449 3019 527 3065
rect 573 3019 651 3065
rect 697 3019 775 3065
rect 821 3019 843 3065
rect 257 2941 843 3019
rect 257 2895 279 2941
rect 325 2895 403 2941
rect 449 2895 527 2941
rect 573 2895 651 2941
rect 697 2895 775 2941
rect 821 2895 843 2941
rect 257 2817 843 2895
rect 257 2771 279 2817
rect 325 2771 403 2817
rect 449 2771 527 2817
rect 573 2771 651 2817
rect 697 2771 775 2817
rect 821 2771 843 2817
rect 257 2693 843 2771
rect 257 2647 279 2693
rect 325 2647 403 2693
rect 449 2647 527 2693
rect 573 2647 651 2693
rect 697 2647 775 2693
rect 821 2647 843 2693
rect 257 2569 843 2647
rect 257 2523 279 2569
rect 325 2523 403 2569
rect 449 2523 527 2569
rect 573 2523 651 2569
rect 697 2523 775 2569
rect 821 2523 843 2569
rect 257 2445 843 2523
rect 257 2399 279 2445
rect 325 2399 403 2445
rect 449 2399 527 2445
rect 573 2399 651 2445
rect 697 2399 775 2445
rect 821 2399 843 2445
rect 257 2321 843 2399
rect 257 2275 279 2321
rect 325 2275 403 2321
rect 449 2275 527 2321
rect 573 2275 651 2321
rect 697 2275 775 2321
rect 821 2275 843 2321
rect 257 2197 843 2275
rect 257 2151 279 2197
rect 325 2151 403 2197
rect 449 2151 527 2197
rect 573 2151 651 2197
rect 697 2151 775 2197
rect 821 2151 843 2197
rect 257 2073 843 2151
rect 257 2027 279 2073
rect 325 2027 403 2073
rect 449 2027 527 2073
rect 573 2027 651 2073
rect 697 2027 775 2073
rect 821 2027 843 2073
rect 257 1949 843 2027
rect 257 1903 279 1949
rect 325 1903 403 1949
rect 449 1903 527 1949
rect 573 1903 651 1949
rect 697 1903 775 1949
rect 821 1903 843 1949
rect 257 1825 843 1903
rect 257 1779 279 1825
rect 325 1779 403 1825
rect 449 1779 527 1825
rect 573 1779 651 1825
rect 697 1779 775 1825
rect 821 1779 843 1825
rect 257 1701 843 1779
rect 257 1655 279 1701
rect 325 1655 403 1701
rect 449 1655 527 1701
rect 573 1655 651 1701
rect 697 1655 775 1701
rect 821 1655 843 1701
rect 257 1577 843 1655
rect 257 1531 279 1577
rect 325 1531 403 1577
rect 449 1531 527 1577
rect 573 1531 651 1577
rect 697 1531 775 1577
rect 821 1531 843 1577
rect 257 1453 843 1531
rect 257 1407 279 1453
rect 325 1407 403 1453
rect 449 1407 527 1453
rect 573 1407 651 1453
rect 697 1407 775 1453
rect 821 1407 843 1453
rect 257 1329 843 1407
rect 257 1283 279 1329
rect 325 1283 403 1329
rect 449 1283 527 1329
rect 573 1283 651 1329
rect 697 1283 775 1329
rect 821 1283 843 1329
rect 257 1205 843 1283
rect 257 1159 279 1205
rect 325 1159 403 1205
rect 449 1159 527 1205
rect 573 1159 651 1205
rect 697 1159 775 1205
rect 821 1159 843 1205
rect 257 1081 843 1159
rect 257 1035 279 1081
rect 325 1035 403 1081
rect 449 1035 527 1081
rect 573 1035 651 1081
rect 697 1035 775 1081
rect 821 1035 843 1081
rect 257 957 843 1035
rect 257 911 279 957
rect 325 911 403 957
rect 449 911 527 957
rect 573 911 651 957
rect 697 911 775 957
rect 821 911 843 957
rect 257 833 843 911
rect 257 787 279 833
rect 325 787 403 833
rect 449 787 527 833
rect 573 787 651 833
rect 697 787 775 833
rect 821 787 843 833
rect 257 709 843 787
rect 257 663 279 709
rect 325 663 403 709
rect 449 663 527 709
rect 573 663 651 709
rect 697 663 775 709
rect 821 663 843 709
rect 257 641 843 663
rect 14203 9265 14939 9287
rect 14203 9219 14225 9265
rect 14271 9219 14349 9265
rect 14395 9219 14473 9265
rect 14519 9219 14597 9265
rect 14643 9219 14721 9265
rect 14767 9219 14939 9265
rect 14203 9141 14939 9219
rect 14203 9095 14225 9141
rect 14271 9095 14349 9141
rect 14395 9095 14473 9141
rect 14519 9095 14597 9141
rect 14643 9095 14721 9141
rect 14767 9095 14939 9141
rect 14203 9017 14939 9095
rect 14203 8971 14225 9017
rect 14271 8971 14349 9017
rect 14395 8971 14473 9017
rect 14519 8971 14597 9017
rect 14643 8971 14721 9017
rect 14767 8971 14939 9017
rect 14203 8893 14939 8971
rect 14203 8847 14225 8893
rect 14271 8847 14349 8893
rect 14395 8847 14473 8893
rect 14519 8847 14597 8893
rect 14643 8847 14721 8893
rect 14767 8847 14939 8893
rect 14203 8769 14939 8847
rect 14203 8723 14225 8769
rect 14271 8723 14349 8769
rect 14395 8723 14473 8769
rect 14519 8723 14597 8769
rect 14643 8723 14721 8769
rect 14767 8723 14939 8769
rect 14203 8645 14939 8723
rect 14203 8599 14225 8645
rect 14271 8599 14349 8645
rect 14395 8599 14473 8645
rect 14519 8599 14597 8645
rect 14643 8599 14721 8645
rect 14767 8599 14939 8645
rect 14203 8521 14939 8599
rect 14203 8475 14225 8521
rect 14271 8475 14349 8521
rect 14395 8475 14473 8521
rect 14519 8475 14597 8521
rect 14643 8475 14721 8521
rect 14767 8475 14939 8521
rect 14203 8397 14939 8475
rect 14203 8351 14225 8397
rect 14271 8351 14349 8397
rect 14395 8351 14473 8397
rect 14519 8351 14597 8397
rect 14643 8351 14721 8397
rect 14767 8351 14939 8397
rect 14203 8273 14939 8351
rect 14203 8227 14225 8273
rect 14271 8227 14349 8273
rect 14395 8227 14473 8273
rect 14519 8227 14597 8273
rect 14643 8227 14721 8273
rect 14767 8227 14939 8273
rect 14203 8149 14939 8227
rect 14203 8103 14225 8149
rect 14271 8103 14349 8149
rect 14395 8103 14473 8149
rect 14519 8103 14597 8149
rect 14643 8103 14721 8149
rect 14767 8103 14939 8149
rect 14203 8025 14939 8103
rect 14203 7979 14225 8025
rect 14271 7979 14349 8025
rect 14395 7979 14473 8025
rect 14519 7979 14597 8025
rect 14643 7979 14721 8025
rect 14767 7979 14939 8025
rect 14203 7901 14939 7979
rect 14203 7855 14225 7901
rect 14271 7855 14349 7901
rect 14395 7855 14473 7901
rect 14519 7855 14597 7901
rect 14643 7855 14721 7901
rect 14767 7855 14939 7901
rect 14203 7777 14939 7855
rect 14203 7731 14225 7777
rect 14271 7731 14349 7777
rect 14395 7731 14473 7777
rect 14519 7731 14597 7777
rect 14643 7731 14721 7777
rect 14767 7731 14939 7777
rect 14203 7653 14939 7731
rect 14203 7607 14225 7653
rect 14271 7607 14349 7653
rect 14395 7607 14473 7653
rect 14519 7607 14597 7653
rect 14643 7607 14721 7653
rect 14767 7607 14939 7653
rect 14203 7529 14939 7607
rect 14203 7483 14225 7529
rect 14271 7483 14349 7529
rect 14395 7483 14473 7529
rect 14519 7483 14597 7529
rect 14643 7483 14721 7529
rect 14767 7483 14939 7529
rect 14203 7405 14939 7483
rect 14203 7359 14225 7405
rect 14271 7359 14349 7405
rect 14395 7359 14473 7405
rect 14519 7359 14597 7405
rect 14643 7359 14721 7405
rect 14767 7359 14939 7405
rect 14203 7281 14939 7359
rect 14203 7235 14225 7281
rect 14271 7235 14349 7281
rect 14395 7235 14473 7281
rect 14519 7235 14597 7281
rect 14643 7235 14721 7281
rect 14767 7235 14939 7281
rect 14203 7157 14939 7235
rect 14203 7111 14225 7157
rect 14271 7111 14349 7157
rect 14395 7111 14473 7157
rect 14519 7111 14597 7157
rect 14643 7111 14721 7157
rect 14767 7111 14939 7157
rect 14203 7033 14939 7111
rect 14203 6987 14225 7033
rect 14271 6987 14349 7033
rect 14395 6987 14473 7033
rect 14519 6987 14597 7033
rect 14643 6987 14721 7033
rect 14767 6987 14939 7033
rect 14203 6909 14939 6987
rect 14203 6863 14225 6909
rect 14271 6863 14349 6909
rect 14395 6863 14473 6909
rect 14519 6863 14597 6909
rect 14643 6863 14721 6909
rect 14767 6863 14939 6909
rect 14203 6785 14939 6863
rect 14203 6739 14225 6785
rect 14271 6739 14349 6785
rect 14395 6739 14473 6785
rect 14519 6739 14597 6785
rect 14643 6739 14721 6785
rect 14767 6739 14939 6785
rect 14203 6661 14939 6739
rect 14203 6615 14225 6661
rect 14271 6615 14349 6661
rect 14395 6615 14473 6661
rect 14519 6615 14597 6661
rect 14643 6615 14721 6661
rect 14767 6615 14939 6661
rect 14203 6537 14939 6615
rect 14203 6491 14225 6537
rect 14271 6491 14349 6537
rect 14395 6491 14473 6537
rect 14519 6491 14597 6537
rect 14643 6491 14721 6537
rect 14767 6491 14939 6537
rect 14203 6413 14939 6491
rect 14203 6367 14225 6413
rect 14271 6367 14349 6413
rect 14395 6367 14473 6413
rect 14519 6367 14597 6413
rect 14643 6367 14721 6413
rect 14767 6367 14939 6413
rect 14203 6289 14939 6367
rect 14203 6243 14225 6289
rect 14271 6243 14349 6289
rect 14395 6243 14473 6289
rect 14519 6243 14597 6289
rect 14643 6243 14721 6289
rect 14767 6243 14939 6289
rect 14203 6165 14939 6243
rect 14203 6119 14225 6165
rect 14271 6119 14349 6165
rect 14395 6119 14473 6165
rect 14519 6119 14597 6165
rect 14643 6119 14721 6165
rect 14767 6119 14939 6165
rect 14203 6041 14939 6119
rect 14203 5995 14225 6041
rect 14271 5995 14349 6041
rect 14395 5995 14473 6041
rect 14519 5995 14597 6041
rect 14643 5995 14721 6041
rect 14767 5995 14939 6041
rect 14203 5917 14939 5995
rect 14203 5871 14225 5917
rect 14271 5871 14349 5917
rect 14395 5871 14473 5917
rect 14519 5871 14597 5917
rect 14643 5871 14721 5917
rect 14767 5871 14939 5917
rect 14203 5793 14939 5871
rect 14203 5747 14225 5793
rect 14271 5747 14349 5793
rect 14395 5747 14473 5793
rect 14519 5747 14597 5793
rect 14643 5747 14721 5793
rect 14767 5747 14939 5793
rect 14203 5669 14939 5747
rect 14203 5623 14225 5669
rect 14271 5623 14349 5669
rect 14395 5623 14473 5669
rect 14519 5623 14597 5669
rect 14643 5623 14721 5669
rect 14767 5623 14939 5669
rect 14203 5545 14939 5623
rect 14203 5499 14225 5545
rect 14271 5499 14349 5545
rect 14395 5499 14473 5545
rect 14519 5499 14597 5545
rect 14643 5499 14721 5545
rect 14767 5499 14939 5545
rect 14203 5421 14939 5499
rect 14203 5375 14225 5421
rect 14271 5375 14349 5421
rect 14395 5375 14473 5421
rect 14519 5375 14597 5421
rect 14643 5375 14721 5421
rect 14767 5375 14939 5421
rect 14203 5297 14939 5375
rect 14203 5251 14225 5297
rect 14271 5251 14349 5297
rect 14395 5251 14473 5297
rect 14519 5251 14597 5297
rect 14643 5251 14721 5297
rect 14767 5251 14939 5297
rect 14203 5173 14939 5251
rect 14203 5127 14225 5173
rect 14271 5127 14349 5173
rect 14395 5127 14473 5173
rect 14519 5127 14597 5173
rect 14643 5127 14721 5173
rect 14767 5127 14939 5173
rect 14203 5049 14939 5127
rect 14203 5003 14225 5049
rect 14271 5003 14349 5049
rect 14395 5003 14473 5049
rect 14519 5003 14597 5049
rect 14643 5003 14721 5049
rect 14767 5003 14939 5049
rect 14203 4925 14939 5003
rect 14203 4879 14225 4925
rect 14271 4879 14349 4925
rect 14395 4879 14473 4925
rect 14519 4879 14597 4925
rect 14643 4879 14721 4925
rect 14767 4879 14939 4925
rect 14203 4801 14939 4879
rect 14203 4755 14225 4801
rect 14271 4755 14349 4801
rect 14395 4755 14473 4801
rect 14519 4755 14597 4801
rect 14643 4755 14721 4801
rect 14767 4755 14939 4801
rect 14203 4677 14939 4755
rect 14203 4631 14225 4677
rect 14271 4631 14349 4677
rect 14395 4631 14473 4677
rect 14519 4631 14597 4677
rect 14643 4631 14721 4677
rect 14767 4631 14939 4677
rect 14203 4553 14939 4631
rect 14203 4507 14225 4553
rect 14271 4507 14349 4553
rect 14395 4507 14473 4553
rect 14519 4507 14597 4553
rect 14643 4507 14721 4553
rect 14767 4507 14939 4553
rect 14203 4429 14939 4507
rect 14203 4383 14225 4429
rect 14271 4383 14349 4429
rect 14395 4383 14473 4429
rect 14519 4383 14597 4429
rect 14643 4383 14721 4429
rect 14767 4383 14939 4429
rect 14203 4305 14939 4383
rect 14203 4259 14225 4305
rect 14271 4259 14349 4305
rect 14395 4259 14473 4305
rect 14519 4259 14597 4305
rect 14643 4259 14721 4305
rect 14767 4259 14939 4305
rect 14203 4181 14939 4259
rect 14203 4135 14225 4181
rect 14271 4135 14349 4181
rect 14395 4135 14473 4181
rect 14519 4135 14597 4181
rect 14643 4135 14721 4181
rect 14767 4135 14939 4181
rect 14203 4057 14939 4135
rect 14203 4011 14225 4057
rect 14271 4011 14349 4057
rect 14395 4011 14473 4057
rect 14519 4011 14597 4057
rect 14643 4011 14721 4057
rect 14767 4011 14939 4057
rect 14203 3933 14939 4011
rect 14203 3887 14225 3933
rect 14271 3887 14349 3933
rect 14395 3887 14473 3933
rect 14519 3887 14597 3933
rect 14643 3887 14721 3933
rect 14767 3887 14939 3933
rect 14203 3809 14939 3887
rect 14203 3763 14225 3809
rect 14271 3763 14349 3809
rect 14395 3763 14473 3809
rect 14519 3763 14597 3809
rect 14643 3763 14721 3809
rect 14767 3763 14939 3809
rect 14203 3685 14939 3763
rect 14203 3639 14225 3685
rect 14271 3639 14349 3685
rect 14395 3639 14473 3685
rect 14519 3639 14597 3685
rect 14643 3639 14721 3685
rect 14767 3639 14939 3685
rect 14203 3561 14939 3639
rect 14203 3515 14225 3561
rect 14271 3515 14349 3561
rect 14395 3515 14473 3561
rect 14519 3515 14597 3561
rect 14643 3515 14721 3561
rect 14767 3515 14939 3561
rect 14203 3437 14939 3515
rect 14203 3391 14225 3437
rect 14271 3391 14349 3437
rect 14395 3391 14473 3437
rect 14519 3391 14597 3437
rect 14643 3391 14721 3437
rect 14767 3391 14939 3437
rect 14203 3313 14939 3391
rect 14203 3267 14225 3313
rect 14271 3267 14349 3313
rect 14395 3267 14473 3313
rect 14519 3267 14597 3313
rect 14643 3267 14721 3313
rect 14767 3267 14939 3313
rect 14203 3189 14939 3267
rect 14203 3143 14225 3189
rect 14271 3143 14349 3189
rect 14395 3143 14473 3189
rect 14519 3143 14597 3189
rect 14643 3143 14721 3189
rect 14767 3143 14939 3189
rect 14203 3065 14939 3143
rect 14203 3019 14225 3065
rect 14271 3019 14349 3065
rect 14395 3019 14473 3065
rect 14519 3019 14597 3065
rect 14643 3019 14721 3065
rect 14767 3019 14939 3065
rect 14203 2941 14939 3019
rect 14203 2895 14225 2941
rect 14271 2895 14349 2941
rect 14395 2895 14473 2941
rect 14519 2895 14597 2941
rect 14643 2895 14721 2941
rect 14767 2895 14939 2941
rect 14203 2817 14939 2895
rect 14203 2771 14225 2817
rect 14271 2771 14349 2817
rect 14395 2771 14473 2817
rect 14519 2771 14597 2817
rect 14643 2771 14721 2817
rect 14767 2771 14939 2817
rect 14203 2693 14939 2771
rect 14203 2647 14225 2693
rect 14271 2647 14349 2693
rect 14395 2647 14473 2693
rect 14519 2647 14597 2693
rect 14643 2647 14721 2693
rect 14767 2647 14939 2693
rect 14203 2569 14939 2647
rect 14203 2523 14225 2569
rect 14271 2523 14349 2569
rect 14395 2523 14473 2569
rect 14519 2523 14597 2569
rect 14643 2523 14721 2569
rect 14767 2523 14939 2569
rect 14203 2445 14939 2523
rect 14203 2399 14225 2445
rect 14271 2399 14349 2445
rect 14395 2399 14473 2445
rect 14519 2399 14597 2445
rect 14643 2399 14721 2445
rect 14767 2399 14939 2445
rect 14203 2321 14939 2399
rect 14203 2275 14225 2321
rect 14271 2275 14349 2321
rect 14395 2275 14473 2321
rect 14519 2275 14597 2321
rect 14643 2275 14721 2321
rect 14767 2275 14939 2321
rect 14203 2197 14939 2275
rect 14203 2151 14225 2197
rect 14271 2151 14349 2197
rect 14395 2151 14473 2197
rect 14519 2151 14597 2197
rect 14643 2151 14721 2197
rect 14767 2151 14939 2197
rect 14203 2073 14939 2151
rect 14203 2027 14225 2073
rect 14271 2027 14349 2073
rect 14395 2027 14473 2073
rect 14519 2027 14597 2073
rect 14643 2027 14721 2073
rect 14767 2027 14939 2073
rect 14203 1949 14939 2027
rect 14203 1903 14225 1949
rect 14271 1903 14349 1949
rect 14395 1903 14473 1949
rect 14519 1903 14597 1949
rect 14643 1903 14721 1949
rect 14767 1903 14939 1949
rect 14203 1825 14939 1903
rect 14203 1779 14225 1825
rect 14271 1779 14349 1825
rect 14395 1779 14473 1825
rect 14519 1779 14597 1825
rect 14643 1779 14721 1825
rect 14767 1779 14939 1825
rect 14203 1701 14939 1779
rect 14203 1655 14225 1701
rect 14271 1655 14349 1701
rect 14395 1655 14473 1701
rect 14519 1655 14597 1701
rect 14643 1655 14721 1701
rect 14767 1655 14939 1701
rect 14203 1577 14939 1655
rect 14203 1531 14225 1577
rect 14271 1531 14349 1577
rect 14395 1531 14473 1577
rect 14519 1531 14597 1577
rect 14643 1531 14721 1577
rect 14767 1531 14939 1577
rect 14203 1453 14939 1531
rect 14203 1407 14225 1453
rect 14271 1407 14349 1453
rect 14395 1407 14473 1453
rect 14519 1407 14597 1453
rect 14643 1407 14721 1453
rect 14767 1407 14939 1453
rect 14203 1329 14939 1407
rect 14203 1283 14225 1329
rect 14271 1283 14349 1329
rect 14395 1283 14473 1329
rect 14519 1283 14597 1329
rect 14643 1283 14721 1329
rect 14767 1283 14939 1329
rect 14203 1205 14939 1283
rect 14203 1159 14225 1205
rect 14271 1159 14349 1205
rect 14395 1159 14473 1205
rect 14519 1159 14597 1205
rect 14643 1159 14721 1205
rect 14767 1159 14939 1205
rect 14203 1081 14939 1159
rect 14203 1035 14225 1081
rect 14271 1035 14349 1081
rect 14395 1035 14473 1081
rect 14519 1035 14597 1081
rect 14643 1035 14721 1081
rect 14767 1035 14939 1081
rect 14203 957 14939 1035
rect 14203 911 14225 957
rect 14271 911 14349 957
rect 14395 911 14473 957
rect 14519 911 14597 957
rect 14643 911 14721 957
rect 14767 911 14939 957
rect 14203 833 14939 911
rect 14203 787 14225 833
rect 14271 787 14349 833
rect 14395 787 14473 833
rect 14519 787 14597 833
rect 14643 787 14721 833
rect 14767 787 14939 833
rect 14203 709 14939 787
rect 14203 663 14225 709
rect 14271 663 14349 709
rect 14395 663 14473 709
rect 14519 663 14597 709
rect 14643 663 14721 709
rect 14767 663 14939 709
rect 14203 641 14939 663
<< nsubdiff >>
rect 1038 55822 2094 55844
rect 1038 54742 1060 55822
rect 1106 55776 1214 55822
rect 1918 55776 2026 55822
rect 1106 55754 2026 55776
rect 1106 54810 1128 55754
rect 2004 54810 2026 55754
rect 1106 54788 2026 54810
rect 1106 54742 1214 54788
rect 1918 54742 2026 54788
rect 2072 54742 2094 55822
rect 1038 54720 2094 54742
<< mvnsubdiff >>
rect 11290 41612 11826 41625
rect 11290 41566 11303 41612
rect 11349 41566 11419 41612
rect 11465 41566 11535 41612
rect 11581 41566 11651 41612
rect 11697 41566 11767 41612
rect 11813 41566 11826 41612
rect 11290 41553 11826 41566
rect 11290 41496 11362 41553
rect 11290 41450 11303 41496
rect 11349 41450 11362 41496
rect 11754 41496 11826 41553
rect 11290 41380 11362 41450
rect 11290 41334 11303 41380
rect 11349 41334 11362 41380
rect 11290 41264 11362 41334
rect 11290 41218 11303 41264
rect 11349 41218 11362 41264
rect 11754 41450 11767 41496
rect 11813 41450 11826 41496
rect 11754 41380 11826 41450
rect 11754 41334 11767 41380
rect 11813 41334 11826 41380
rect 11754 41264 11826 41334
rect 11290 41161 11362 41218
rect 11754 41218 11767 41264
rect 11813 41218 11826 41264
rect 11754 41161 11826 41218
rect 11290 41148 11826 41161
rect 11290 41102 11303 41148
rect 11349 41102 11419 41148
rect 11465 41102 11535 41148
rect 11581 41102 11651 41148
rect 11697 41102 11767 41148
rect 11813 41102 11826 41148
rect 11290 41089 11826 41102
rect 11290 41032 11362 41089
rect 11290 40986 11303 41032
rect 11349 40986 11362 41032
rect 11754 41032 11826 41089
rect 11290 40916 11362 40986
rect 11290 40870 11303 40916
rect 11349 40870 11362 40916
rect 11290 40800 11362 40870
rect 11290 40754 11303 40800
rect 11349 40754 11362 40800
rect 11754 40986 11767 41032
rect 11813 40986 11826 41032
rect 11754 40916 11826 40986
rect 11754 40870 11767 40916
rect 11813 40870 11826 40916
rect 11754 40800 11826 40870
rect 11290 40697 11362 40754
rect 11754 40754 11767 40800
rect 11813 40754 11826 40800
rect 11754 40697 11826 40754
rect 11290 40684 11826 40697
rect 11290 40638 11303 40684
rect 11349 40638 11419 40684
rect 11465 40638 11535 40684
rect 11581 40638 11651 40684
rect 11697 40638 11767 40684
rect 11813 40638 11826 40684
rect 11290 40625 11826 40638
<< psubdiffcont >>
rect 2353 56786 14713 56832
rect 2353 55870 2399 56668
rect 14667 55870 14713 56668
rect 2353 55706 14713 55752
rect 10764 43212 10810 43258
rect 10878 43212 10924 43258
rect 10992 43212 11038 43258
rect 11106 43212 11152 43258
rect 11220 43212 11266 43258
rect 11334 43212 11380 43258
rect 11448 43212 11494 43258
rect 11562 43212 11608 43258
rect 11676 43212 11722 43258
rect 11790 43212 11836 43258
rect 10764 43098 10810 43144
rect 10878 43098 10924 43144
rect 10992 43098 11038 43144
rect 11106 43098 11152 43144
rect 11220 43098 11266 43144
rect 11334 43098 11380 43144
rect 11448 43098 11494 43144
rect 11562 43098 11608 43144
rect 11676 43098 11722 43144
rect 11790 43098 11836 43144
rect 10764 42984 10810 43030
rect 10878 42984 10924 43030
rect 10992 42984 11038 43030
rect 11106 42984 11152 43030
rect 11220 42984 11266 43030
rect 11334 42984 11380 43030
rect 11448 42984 11494 43030
rect 11562 42984 11608 43030
rect 11676 42984 11722 43030
rect 11790 42984 11836 43030
rect 10764 42870 10810 42916
rect 10878 42870 10924 42916
rect 10992 42870 11038 42916
rect 11106 42870 11152 42916
rect 11220 42870 11266 42916
rect 11334 42870 11380 42916
rect 11448 42870 11494 42916
rect 11562 42870 11608 42916
rect 11676 42870 11722 42916
rect 11790 42870 11836 42916
rect 10764 42756 10810 42802
rect 10878 42756 10924 42802
rect 10992 42756 11038 42802
rect 11106 42756 11152 42802
rect 11220 42756 11266 42802
rect 11334 42756 11380 42802
rect 11448 42756 11494 42802
rect 11562 42756 11608 42802
rect 11676 42756 11722 42802
rect 11790 42756 11836 42802
rect 10764 42642 10810 42688
rect 10878 42642 10924 42688
rect 10992 42642 11038 42688
rect 11106 42642 11152 42688
rect 11220 42642 11266 42688
rect 11334 42642 11380 42688
rect 11448 42642 11494 42688
rect 11562 42642 11608 42688
rect 11676 42642 11722 42688
rect 11790 42642 11836 42688
rect 10764 42528 10810 42574
rect 10878 42528 10924 42574
rect 10992 42528 11038 42574
rect 11106 42528 11152 42574
rect 11220 42528 11266 42574
rect 11334 42528 11380 42574
rect 11448 42528 11494 42574
rect 11562 42528 11608 42574
rect 11676 42528 11722 42574
rect 11790 42528 11836 42574
rect 10764 42414 10810 42460
rect 10878 42414 10924 42460
rect 10992 42414 11038 42460
rect 11106 42414 11152 42460
rect 11220 42414 11266 42460
rect 11334 42414 11380 42460
rect 11448 42414 11494 42460
rect 11562 42414 11608 42460
rect 11676 42414 11722 42460
rect 11790 42414 11836 42460
rect 10764 42300 10810 42346
rect 10878 42300 10924 42346
rect 10992 42300 11038 42346
rect 11106 42300 11152 42346
rect 11220 42300 11266 42346
rect 11334 42300 11380 42346
rect 11448 42300 11494 42346
rect 11562 42300 11608 42346
rect 11676 42300 11722 42346
rect 11790 42300 11836 42346
rect 12075 40717 12121 43207
rect 12182 43161 14484 43207
rect 12182 40717 14484 40763
rect 14592 40717 14638 43207
rect 279 9219 325 9265
rect 403 9219 449 9265
rect 527 9219 573 9265
rect 651 9219 697 9265
rect 775 9219 821 9265
rect 279 9095 325 9141
rect 403 9095 449 9141
rect 527 9095 573 9141
rect 651 9095 697 9141
rect 775 9095 821 9141
rect 279 8971 325 9017
rect 403 8971 449 9017
rect 527 8971 573 9017
rect 651 8971 697 9017
rect 775 8971 821 9017
rect 279 8847 325 8893
rect 403 8847 449 8893
rect 527 8847 573 8893
rect 651 8847 697 8893
rect 775 8847 821 8893
rect 279 8723 325 8769
rect 403 8723 449 8769
rect 527 8723 573 8769
rect 651 8723 697 8769
rect 775 8723 821 8769
rect 279 8599 325 8645
rect 403 8599 449 8645
rect 527 8599 573 8645
rect 651 8599 697 8645
rect 775 8599 821 8645
rect 279 8475 325 8521
rect 403 8475 449 8521
rect 527 8475 573 8521
rect 651 8475 697 8521
rect 775 8475 821 8521
rect 279 8351 325 8397
rect 403 8351 449 8397
rect 527 8351 573 8397
rect 651 8351 697 8397
rect 775 8351 821 8397
rect 279 8227 325 8273
rect 403 8227 449 8273
rect 527 8227 573 8273
rect 651 8227 697 8273
rect 775 8227 821 8273
rect 279 8103 325 8149
rect 403 8103 449 8149
rect 527 8103 573 8149
rect 651 8103 697 8149
rect 775 8103 821 8149
rect 279 7979 325 8025
rect 403 7979 449 8025
rect 527 7979 573 8025
rect 651 7979 697 8025
rect 775 7979 821 8025
rect 279 7855 325 7901
rect 403 7855 449 7901
rect 527 7855 573 7901
rect 651 7855 697 7901
rect 775 7855 821 7901
rect 279 7731 325 7777
rect 403 7731 449 7777
rect 527 7731 573 7777
rect 651 7731 697 7777
rect 775 7731 821 7777
rect 279 7607 325 7653
rect 403 7607 449 7653
rect 527 7607 573 7653
rect 651 7607 697 7653
rect 775 7607 821 7653
rect 279 7483 325 7529
rect 403 7483 449 7529
rect 527 7483 573 7529
rect 651 7483 697 7529
rect 775 7483 821 7529
rect 279 7359 325 7405
rect 403 7359 449 7405
rect 527 7359 573 7405
rect 651 7359 697 7405
rect 775 7359 821 7405
rect 279 7235 325 7281
rect 403 7235 449 7281
rect 527 7235 573 7281
rect 651 7235 697 7281
rect 775 7235 821 7281
rect 279 7111 325 7157
rect 403 7111 449 7157
rect 527 7111 573 7157
rect 651 7111 697 7157
rect 775 7111 821 7157
rect 279 6987 325 7033
rect 403 6987 449 7033
rect 527 6987 573 7033
rect 651 6987 697 7033
rect 775 6987 821 7033
rect 279 6863 325 6909
rect 403 6863 449 6909
rect 527 6863 573 6909
rect 651 6863 697 6909
rect 775 6863 821 6909
rect 279 6739 325 6785
rect 403 6739 449 6785
rect 527 6739 573 6785
rect 651 6739 697 6785
rect 775 6739 821 6785
rect 279 6615 325 6661
rect 403 6615 449 6661
rect 527 6615 573 6661
rect 651 6615 697 6661
rect 775 6615 821 6661
rect 279 6491 325 6537
rect 403 6491 449 6537
rect 527 6491 573 6537
rect 651 6491 697 6537
rect 775 6491 821 6537
rect 279 6367 325 6413
rect 403 6367 449 6413
rect 527 6367 573 6413
rect 651 6367 697 6413
rect 775 6367 821 6413
rect 279 6243 325 6289
rect 403 6243 449 6289
rect 527 6243 573 6289
rect 651 6243 697 6289
rect 775 6243 821 6289
rect 279 6119 325 6165
rect 403 6119 449 6165
rect 527 6119 573 6165
rect 651 6119 697 6165
rect 775 6119 821 6165
rect 279 5995 325 6041
rect 403 5995 449 6041
rect 527 5995 573 6041
rect 651 5995 697 6041
rect 775 5995 821 6041
rect 279 5871 325 5917
rect 403 5871 449 5917
rect 527 5871 573 5917
rect 651 5871 697 5917
rect 775 5871 821 5917
rect 279 5747 325 5793
rect 403 5747 449 5793
rect 527 5747 573 5793
rect 651 5747 697 5793
rect 775 5747 821 5793
rect 279 5623 325 5669
rect 403 5623 449 5669
rect 527 5623 573 5669
rect 651 5623 697 5669
rect 775 5623 821 5669
rect 279 5499 325 5545
rect 403 5499 449 5545
rect 527 5499 573 5545
rect 651 5499 697 5545
rect 775 5499 821 5545
rect 279 5375 325 5421
rect 403 5375 449 5421
rect 527 5375 573 5421
rect 651 5375 697 5421
rect 775 5375 821 5421
rect 279 5251 325 5297
rect 403 5251 449 5297
rect 527 5251 573 5297
rect 651 5251 697 5297
rect 775 5251 821 5297
rect 279 5127 325 5173
rect 403 5127 449 5173
rect 527 5127 573 5173
rect 651 5127 697 5173
rect 775 5127 821 5173
rect 279 5003 325 5049
rect 403 5003 449 5049
rect 527 5003 573 5049
rect 651 5003 697 5049
rect 775 5003 821 5049
rect 279 4879 325 4925
rect 403 4879 449 4925
rect 527 4879 573 4925
rect 651 4879 697 4925
rect 775 4879 821 4925
rect 279 4755 325 4801
rect 403 4755 449 4801
rect 527 4755 573 4801
rect 651 4755 697 4801
rect 775 4755 821 4801
rect 279 4631 325 4677
rect 403 4631 449 4677
rect 527 4631 573 4677
rect 651 4631 697 4677
rect 775 4631 821 4677
rect 279 4507 325 4553
rect 403 4507 449 4553
rect 527 4507 573 4553
rect 651 4507 697 4553
rect 775 4507 821 4553
rect 279 4383 325 4429
rect 403 4383 449 4429
rect 527 4383 573 4429
rect 651 4383 697 4429
rect 775 4383 821 4429
rect 279 4259 325 4305
rect 403 4259 449 4305
rect 527 4259 573 4305
rect 651 4259 697 4305
rect 775 4259 821 4305
rect 279 4135 325 4181
rect 403 4135 449 4181
rect 527 4135 573 4181
rect 651 4135 697 4181
rect 775 4135 821 4181
rect 279 4011 325 4057
rect 403 4011 449 4057
rect 527 4011 573 4057
rect 651 4011 697 4057
rect 775 4011 821 4057
rect 279 3887 325 3933
rect 403 3887 449 3933
rect 527 3887 573 3933
rect 651 3887 697 3933
rect 775 3887 821 3933
rect 279 3763 325 3809
rect 403 3763 449 3809
rect 527 3763 573 3809
rect 651 3763 697 3809
rect 775 3763 821 3809
rect 279 3639 325 3685
rect 403 3639 449 3685
rect 527 3639 573 3685
rect 651 3639 697 3685
rect 775 3639 821 3685
rect 279 3515 325 3561
rect 403 3515 449 3561
rect 527 3515 573 3561
rect 651 3515 697 3561
rect 775 3515 821 3561
rect 279 3391 325 3437
rect 403 3391 449 3437
rect 527 3391 573 3437
rect 651 3391 697 3437
rect 775 3391 821 3437
rect 279 3267 325 3313
rect 403 3267 449 3313
rect 527 3267 573 3313
rect 651 3267 697 3313
rect 775 3267 821 3313
rect 279 3143 325 3189
rect 403 3143 449 3189
rect 527 3143 573 3189
rect 651 3143 697 3189
rect 775 3143 821 3189
rect 279 3019 325 3065
rect 403 3019 449 3065
rect 527 3019 573 3065
rect 651 3019 697 3065
rect 775 3019 821 3065
rect 279 2895 325 2941
rect 403 2895 449 2941
rect 527 2895 573 2941
rect 651 2895 697 2941
rect 775 2895 821 2941
rect 279 2771 325 2817
rect 403 2771 449 2817
rect 527 2771 573 2817
rect 651 2771 697 2817
rect 775 2771 821 2817
rect 279 2647 325 2693
rect 403 2647 449 2693
rect 527 2647 573 2693
rect 651 2647 697 2693
rect 775 2647 821 2693
rect 279 2523 325 2569
rect 403 2523 449 2569
rect 527 2523 573 2569
rect 651 2523 697 2569
rect 775 2523 821 2569
rect 279 2399 325 2445
rect 403 2399 449 2445
rect 527 2399 573 2445
rect 651 2399 697 2445
rect 775 2399 821 2445
rect 279 2275 325 2321
rect 403 2275 449 2321
rect 527 2275 573 2321
rect 651 2275 697 2321
rect 775 2275 821 2321
rect 279 2151 325 2197
rect 403 2151 449 2197
rect 527 2151 573 2197
rect 651 2151 697 2197
rect 775 2151 821 2197
rect 279 2027 325 2073
rect 403 2027 449 2073
rect 527 2027 573 2073
rect 651 2027 697 2073
rect 775 2027 821 2073
rect 279 1903 325 1949
rect 403 1903 449 1949
rect 527 1903 573 1949
rect 651 1903 697 1949
rect 775 1903 821 1949
rect 279 1779 325 1825
rect 403 1779 449 1825
rect 527 1779 573 1825
rect 651 1779 697 1825
rect 775 1779 821 1825
rect 279 1655 325 1701
rect 403 1655 449 1701
rect 527 1655 573 1701
rect 651 1655 697 1701
rect 775 1655 821 1701
rect 279 1531 325 1577
rect 403 1531 449 1577
rect 527 1531 573 1577
rect 651 1531 697 1577
rect 775 1531 821 1577
rect 279 1407 325 1453
rect 403 1407 449 1453
rect 527 1407 573 1453
rect 651 1407 697 1453
rect 775 1407 821 1453
rect 279 1283 325 1329
rect 403 1283 449 1329
rect 527 1283 573 1329
rect 651 1283 697 1329
rect 775 1283 821 1329
rect 279 1159 325 1205
rect 403 1159 449 1205
rect 527 1159 573 1205
rect 651 1159 697 1205
rect 775 1159 821 1205
rect 279 1035 325 1081
rect 403 1035 449 1081
rect 527 1035 573 1081
rect 651 1035 697 1081
rect 775 1035 821 1081
rect 279 911 325 957
rect 403 911 449 957
rect 527 911 573 957
rect 651 911 697 957
rect 775 911 821 957
rect 279 787 325 833
rect 403 787 449 833
rect 527 787 573 833
rect 651 787 697 833
rect 775 787 821 833
rect 279 663 325 709
rect 403 663 449 709
rect 527 663 573 709
rect 651 663 697 709
rect 775 663 821 709
rect 14225 9219 14271 9265
rect 14349 9219 14395 9265
rect 14473 9219 14519 9265
rect 14597 9219 14643 9265
rect 14721 9219 14767 9265
rect 14225 9095 14271 9141
rect 14349 9095 14395 9141
rect 14473 9095 14519 9141
rect 14597 9095 14643 9141
rect 14721 9095 14767 9141
rect 14225 8971 14271 9017
rect 14349 8971 14395 9017
rect 14473 8971 14519 9017
rect 14597 8971 14643 9017
rect 14721 8971 14767 9017
rect 14225 8847 14271 8893
rect 14349 8847 14395 8893
rect 14473 8847 14519 8893
rect 14597 8847 14643 8893
rect 14721 8847 14767 8893
rect 14225 8723 14271 8769
rect 14349 8723 14395 8769
rect 14473 8723 14519 8769
rect 14597 8723 14643 8769
rect 14721 8723 14767 8769
rect 14225 8599 14271 8645
rect 14349 8599 14395 8645
rect 14473 8599 14519 8645
rect 14597 8599 14643 8645
rect 14721 8599 14767 8645
rect 14225 8475 14271 8521
rect 14349 8475 14395 8521
rect 14473 8475 14519 8521
rect 14597 8475 14643 8521
rect 14721 8475 14767 8521
rect 14225 8351 14271 8397
rect 14349 8351 14395 8397
rect 14473 8351 14519 8397
rect 14597 8351 14643 8397
rect 14721 8351 14767 8397
rect 14225 8227 14271 8273
rect 14349 8227 14395 8273
rect 14473 8227 14519 8273
rect 14597 8227 14643 8273
rect 14721 8227 14767 8273
rect 14225 8103 14271 8149
rect 14349 8103 14395 8149
rect 14473 8103 14519 8149
rect 14597 8103 14643 8149
rect 14721 8103 14767 8149
rect 14225 7979 14271 8025
rect 14349 7979 14395 8025
rect 14473 7979 14519 8025
rect 14597 7979 14643 8025
rect 14721 7979 14767 8025
rect 14225 7855 14271 7901
rect 14349 7855 14395 7901
rect 14473 7855 14519 7901
rect 14597 7855 14643 7901
rect 14721 7855 14767 7901
rect 14225 7731 14271 7777
rect 14349 7731 14395 7777
rect 14473 7731 14519 7777
rect 14597 7731 14643 7777
rect 14721 7731 14767 7777
rect 14225 7607 14271 7653
rect 14349 7607 14395 7653
rect 14473 7607 14519 7653
rect 14597 7607 14643 7653
rect 14721 7607 14767 7653
rect 14225 7483 14271 7529
rect 14349 7483 14395 7529
rect 14473 7483 14519 7529
rect 14597 7483 14643 7529
rect 14721 7483 14767 7529
rect 14225 7359 14271 7405
rect 14349 7359 14395 7405
rect 14473 7359 14519 7405
rect 14597 7359 14643 7405
rect 14721 7359 14767 7405
rect 14225 7235 14271 7281
rect 14349 7235 14395 7281
rect 14473 7235 14519 7281
rect 14597 7235 14643 7281
rect 14721 7235 14767 7281
rect 14225 7111 14271 7157
rect 14349 7111 14395 7157
rect 14473 7111 14519 7157
rect 14597 7111 14643 7157
rect 14721 7111 14767 7157
rect 14225 6987 14271 7033
rect 14349 6987 14395 7033
rect 14473 6987 14519 7033
rect 14597 6987 14643 7033
rect 14721 6987 14767 7033
rect 14225 6863 14271 6909
rect 14349 6863 14395 6909
rect 14473 6863 14519 6909
rect 14597 6863 14643 6909
rect 14721 6863 14767 6909
rect 14225 6739 14271 6785
rect 14349 6739 14395 6785
rect 14473 6739 14519 6785
rect 14597 6739 14643 6785
rect 14721 6739 14767 6785
rect 14225 6615 14271 6661
rect 14349 6615 14395 6661
rect 14473 6615 14519 6661
rect 14597 6615 14643 6661
rect 14721 6615 14767 6661
rect 14225 6491 14271 6537
rect 14349 6491 14395 6537
rect 14473 6491 14519 6537
rect 14597 6491 14643 6537
rect 14721 6491 14767 6537
rect 14225 6367 14271 6413
rect 14349 6367 14395 6413
rect 14473 6367 14519 6413
rect 14597 6367 14643 6413
rect 14721 6367 14767 6413
rect 14225 6243 14271 6289
rect 14349 6243 14395 6289
rect 14473 6243 14519 6289
rect 14597 6243 14643 6289
rect 14721 6243 14767 6289
rect 14225 6119 14271 6165
rect 14349 6119 14395 6165
rect 14473 6119 14519 6165
rect 14597 6119 14643 6165
rect 14721 6119 14767 6165
rect 14225 5995 14271 6041
rect 14349 5995 14395 6041
rect 14473 5995 14519 6041
rect 14597 5995 14643 6041
rect 14721 5995 14767 6041
rect 14225 5871 14271 5917
rect 14349 5871 14395 5917
rect 14473 5871 14519 5917
rect 14597 5871 14643 5917
rect 14721 5871 14767 5917
rect 14225 5747 14271 5793
rect 14349 5747 14395 5793
rect 14473 5747 14519 5793
rect 14597 5747 14643 5793
rect 14721 5747 14767 5793
rect 14225 5623 14271 5669
rect 14349 5623 14395 5669
rect 14473 5623 14519 5669
rect 14597 5623 14643 5669
rect 14721 5623 14767 5669
rect 14225 5499 14271 5545
rect 14349 5499 14395 5545
rect 14473 5499 14519 5545
rect 14597 5499 14643 5545
rect 14721 5499 14767 5545
rect 14225 5375 14271 5421
rect 14349 5375 14395 5421
rect 14473 5375 14519 5421
rect 14597 5375 14643 5421
rect 14721 5375 14767 5421
rect 14225 5251 14271 5297
rect 14349 5251 14395 5297
rect 14473 5251 14519 5297
rect 14597 5251 14643 5297
rect 14721 5251 14767 5297
rect 14225 5127 14271 5173
rect 14349 5127 14395 5173
rect 14473 5127 14519 5173
rect 14597 5127 14643 5173
rect 14721 5127 14767 5173
rect 14225 5003 14271 5049
rect 14349 5003 14395 5049
rect 14473 5003 14519 5049
rect 14597 5003 14643 5049
rect 14721 5003 14767 5049
rect 14225 4879 14271 4925
rect 14349 4879 14395 4925
rect 14473 4879 14519 4925
rect 14597 4879 14643 4925
rect 14721 4879 14767 4925
rect 14225 4755 14271 4801
rect 14349 4755 14395 4801
rect 14473 4755 14519 4801
rect 14597 4755 14643 4801
rect 14721 4755 14767 4801
rect 14225 4631 14271 4677
rect 14349 4631 14395 4677
rect 14473 4631 14519 4677
rect 14597 4631 14643 4677
rect 14721 4631 14767 4677
rect 14225 4507 14271 4553
rect 14349 4507 14395 4553
rect 14473 4507 14519 4553
rect 14597 4507 14643 4553
rect 14721 4507 14767 4553
rect 14225 4383 14271 4429
rect 14349 4383 14395 4429
rect 14473 4383 14519 4429
rect 14597 4383 14643 4429
rect 14721 4383 14767 4429
rect 14225 4259 14271 4305
rect 14349 4259 14395 4305
rect 14473 4259 14519 4305
rect 14597 4259 14643 4305
rect 14721 4259 14767 4305
rect 14225 4135 14271 4181
rect 14349 4135 14395 4181
rect 14473 4135 14519 4181
rect 14597 4135 14643 4181
rect 14721 4135 14767 4181
rect 14225 4011 14271 4057
rect 14349 4011 14395 4057
rect 14473 4011 14519 4057
rect 14597 4011 14643 4057
rect 14721 4011 14767 4057
rect 14225 3887 14271 3933
rect 14349 3887 14395 3933
rect 14473 3887 14519 3933
rect 14597 3887 14643 3933
rect 14721 3887 14767 3933
rect 14225 3763 14271 3809
rect 14349 3763 14395 3809
rect 14473 3763 14519 3809
rect 14597 3763 14643 3809
rect 14721 3763 14767 3809
rect 14225 3639 14271 3685
rect 14349 3639 14395 3685
rect 14473 3639 14519 3685
rect 14597 3639 14643 3685
rect 14721 3639 14767 3685
rect 14225 3515 14271 3561
rect 14349 3515 14395 3561
rect 14473 3515 14519 3561
rect 14597 3515 14643 3561
rect 14721 3515 14767 3561
rect 14225 3391 14271 3437
rect 14349 3391 14395 3437
rect 14473 3391 14519 3437
rect 14597 3391 14643 3437
rect 14721 3391 14767 3437
rect 14225 3267 14271 3313
rect 14349 3267 14395 3313
rect 14473 3267 14519 3313
rect 14597 3267 14643 3313
rect 14721 3267 14767 3313
rect 14225 3143 14271 3189
rect 14349 3143 14395 3189
rect 14473 3143 14519 3189
rect 14597 3143 14643 3189
rect 14721 3143 14767 3189
rect 14225 3019 14271 3065
rect 14349 3019 14395 3065
rect 14473 3019 14519 3065
rect 14597 3019 14643 3065
rect 14721 3019 14767 3065
rect 14225 2895 14271 2941
rect 14349 2895 14395 2941
rect 14473 2895 14519 2941
rect 14597 2895 14643 2941
rect 14721 2895 14767 2941
rect 14225 2771 14271 2817
rect 14349 2771 14395 2817
rect 14473 2771 14519 2817
rect 14597 2771 14643 2817
rect 14721 2771 14767 2817
rect 14225 2647 14271 2693
rect 14349 2647 14395 2693
rect 14473 2647 14519 2693
rect 14597 2647 14643 2693
rect 14721 2647 14767 2693
rect 14225 2523 14271 2569
rect 14349 2523 14395 2569
rect 14473 2523 14519 2569
rect 14597 2523 14643 2569
rect 14721 2523 14767 2569
rect 14225 2399 14271 2445
rect 14349 2399 14395 2445
rect 14473 2399 14519 2445
rect 14597 2399 14643 2445
rect 14721 2399 14767 2445
rect 14225 2275 14271 2321
rect 14349 2275 14395 2321
rect 14473 2275 14519 2321
rect 14597 2275 14643 2321
rect 14721 2275 14767 2321
rect 14225 2151 14271 2197
rect 14349 2151 14395 2197
rect 14473 2151 14519 2197
rect 14597 2151 14643 2197
rect 14721 2151 14767 2197
rect 14225 2027 14271 2073
rect 14349 2027 14395 2073
rect 14473 2027 14519 2073
rect 14597 2027 14643 2073
rect 14721 2027 14767 2073
rect 14225 1903 14271 1949
rect 14349 1903 14395 1949
rect 14473 1903 14519 1949
rect 14597 1903 14643 1949
rect 14721 1903 14767 1949
rect 14225 1779 14271 1825
rect 14349 1779 14395 1825
rect 14473 1779 14519 1825
rect 14597 1779 14643 1825
rect 14721 1779 14767 1825
rect 14225 1655 14271 1701
rect 14349 1655 14395 1701
rect 14473 1655 14519 1701
rect 14597 1655 14643 1701
rect 14721 1655 14767 1701
rect 14225 1531 14271 1577
rect 14349 1531 14395 1577
rect 14473 1531 14519 1577
rect 14597 1531 14643 1577
rect 14721 1531 14767 1577
rect 14225 1407 14271 1453
rect 14349 1407 14395 1453
rect 14473 1407 14519 1453
rect 14597 1407 14643 1453
rect 14721 1407 14767 1453
rect 14225 1283 14271 1329
rect 14349 1283 14395 1329
rect 14473 1283 14519 1329
rect 14597 1283 14643 1329
rect 14721 1283 14767 1329
rect 14225 1159 14271 1205
rect 14349 1159 14395 1205
rect 14473 1159 14519 1205
rect 14597 1159 14643 1205
rect 14721 1159 14767 1205
rect 14225 1035 14271 1081
rect 14349 1035 14395 1081
rect 14473 1035 14519 1081
rect 14597 1035 14643 1081
rect 14721 1035 14767 1081
rect 14225 911 14271 957
rect 14349 911 14395 957
rect 14473 911 14519 957
rect 14597 911 14643 957
rect 14721 911 14767 957
rect 14225 787 14271 833
rect 14349 787 14395 833
rect 14473 787 14519 833
rect 14597 787 14643 833
rect 14721 787 14767 833
rect 14225 663 14271 709
rect 14349 663 14395 709
rect 14473 663 14519 709
rect 14597 663 14643 709
rect 14721 663 14767 709
<< nsubdiffcont >>
rect 1060 54742 1106 55822
rect 1214 55776 1918 55822
rect 1214 54742 1918 54788
rect 2026 54742 2072 55822
<< mvnsubdiffcont >>
rect 11303 41566 11349 41612
rect 11419 41566 11465 41612
rect 11535 41566 11581 41612
rect 11651 41566 11697 41612
rect 11767 41566 11813 41612
rect 11303 41450 11349 41496
rect 11303 41334 11349 41380
rect 11303 41218 11349 41264
rect 11767 41450 11813 41496
rect 11767 41334 11813 41380
rect 11767 41218 11813 41264
rect 11303 41102 11349 41148
rect 11419 41102 11465 41148
rect 11535 41102 11581 41148
rect 11651 41102 11697 41148
rect 11767 41102 11813 41148
rect 11303 40986 11349 41032
rect 11303 40870 11349 40916
rect 11303 40754 11349 40800
rect 11767 40986 11813 41032
rect 11767 40870 11813 40916
rect 11767 40754 11813 40800
rect 11303 40638 11349 40684
rect 11419 40638 11465 40684
rect 11535 40638 11581 40684
rect 11651 40638 11697 40684
rect 11767 40638 11813 40684
<< mvnmoscap >>
rect 2760 56119 3760 56419
rect 4260 56119 5260 56419
rect 5760 56119 6760 56419
rect 7260 56119 8260 56419
rect 8760 56119 9760 56419
rect 10260 56119 11260 56419
rect 11760 56119 12760 56419
rect 13260 56119 14260 56419
rect 12482 42146 13082 42746
rect 13622 42146 14222 42746
rect 12482 41178 13082 41778
rect 13622 41178 14222 41778
<< polysilicon >>
rect 2668 56366 2760 56419
rect 2668 56320 2681 56366
rect 2727 56320 2760 56366
rect 2668 56218 2760 56320
rect 2668 56172 2681 56218
rect 2727 56172 2760 56218
rect 2668 56119 2760 56172
rect 3760 56366 3852 56419
rect 3760 56320 3793 56366
rect 3839 56320 3852 56366
rect 3760 56218 3852 56320
rect 3760 56172 3793 56218
rect 3839 56172 3852 56218
rect 3760 56119 3852 56172
rect 4168 56366 4260 56419
rect 4168 56320 4181 56366
rect 4227 56320 4260 56366
rect 4168 56218 4260 56320
rect 4168 56172 4181 56218
rect 4227 56172 4260 56218
rect 4168 56119 4260 56172
rect 5260 56366 5352 56419
rect 5260 56320 5293 56366
rect 5339 56320 5352 56366
rect 5260 56218 5352 56320
rect 5260 56172 5293 56218
rect 5339 56172 5352 56218
rect 5260 56119 5352 56172
rect 5668 56366 5760 56419
rect 5668 56320 5681 56366
rect 5727 56320 5760 56366
rect 5668 56218 5760 56320
rect 5668 56172 5681 56218
rect 5727 56172 5760 56218
rect 5668 56119 5760 56172
rect 6760 56366 6852 56419
rect 6760 56320 6793 56366
rect 6839 56320 6852 56366
rect 6760 56218 6852 56320
rect 6760 56172 6793 56218
rect 6839 56172 6852 56218
rect 6760 56119 6852 56172
rect 7168 56366 7260 56419
rect 7168 56320 7181 56366
rect 7227 56320 7260 56366
rect 7168 56218 7260 56320
rect 7168 56172 7181 56218
rect 7227 56172 7260 56218
rect 7168 56119 7260 56172
rect 8260 56366 8352 56419
rect 8260 56320 8293 56366
rect 8339 56320 8352 56366
rect 8260 56218 8352 56320
rect 8260 56172 8293 56218
rect 8339 56172 8352 56218
rect 8260 56119 8352 56172
rect 8668 56366 8760 56419
rect 8668 56320 8681 56366
rect 8727 56320 8760 56366
rect 8668 56218 8760 56320
rect 8668 56172 8681 56218
rect 8727 56172 8760 56218
rect 8668 56119 8760 56172
rect 9760 56366 9852 56419
rect 9760 56320 9793 56366
rect 9839 56320 9852 56366
rect 9760 56218 9852 56320
rect 9760 56172 9793 56218
rect 9839 56172 9852 56218
rect 9760 56119 9852 56172
rect 10168 56366 10260 56419
rect 10168 56320 10181 56366
rect 10227 56320 10260 56366
rect 10168 56218 10260 56320
rect 10168 56172 10181 56218
rect 10227 56172 10260 56218
rect 10168 56119 10260 56172
rect 11260 56366 11352 56419
rect 11260 56320 11293 56366
rect 11339 56320 11352 56366
rect 11260 56218 11352 56320
rect 11260 56172 11293 56218
rect 11339 56172 11352 56218
rect 11260 56119 11352 56172
rect 11668 56366 11760 56419
rect 11668 56320 11681 56366
rect 11727 56320 11760 56366
rect 11668 56218 11760 56320
rect 11668 56172 11681 56218
rect 11727 56172 11760 56218
rect 11668 56119 11760 56172
rect 12760 56366 12852 56419
rect 12760 56320 12793 56366
rect 12839 56320 12852 56366
rect 12760 56218 12852 56320
rect 12760 56172 12793 56218
rect 12839 56172 12852 56218
rect 12760 56119 12852 56172
rect 13168 56366 13260 56419
rect 13168 56320 13181 56366
rect 13227 56320 13260 56366
rect 13168 56218 13260 56320
rect 13168 56172 13181 56218
rect 13227 56172 13260 56218
rect 13168 56119 13260 56172
rect 14260 56366 14352 56419
rect 14260 56320 14293 56366
rect 14339 56320 14352 56366
rect 14260 56218 14352 56320
rect 14260 56172 14293 56218
rect 14339 56172 14352 56218
rect 14260 56119 14352 56172
rect 1346 55531 1506 55544
rect 1346 55485 1403 55531
rect 1449 55485 1506 55531
rect 1346 55442 1506 55485
rect 1346 55079 1506 55122
rect 1346 55033 1403 55079
rect 1449 55033 1506 55079
rect 1346 55020 1506 55033
rect 1626 55531 1786 55544
rect 1626 55485 1683 55531
rect 1729 55485 1786 55531
rect 1626 55442 1786 55485
rect 1626 55079 1786 55122
rect 1626 55033 1683 55079
rect 1729 55033 1786 55079
rect 1626 55020 1786 55033
rect 12390 42693 12482 42746
rect 12390 42647 12403 42693
rect 12449 42647 12482 42693
rect 12390 42581 12482 42647
rect 12390 42535 12403 42581
rect 12449 42535 12482 42581
rect 12390 42469 12482 42535
rect 12390 42423 12403 42469
rect 12449 42423 12482 42469
rect 12390 42357 12482 42423
rect 12390 42311 12403 42357
rect 12449 42311 12482 42357
rect 12390 42245 12482 42311
rect 12390 42199 12403 42245
rect 12449 42199 12482 42245
rect 12390 42146 12482 42199
rect 13082 42693 13174 42746
rect 13082 42647 13115 42693
rect 13161 42647 13174 42693
rect 13082 42581 13174 42647
rect 13082 42535 13115 42581
rect 13161 42535 13174 42581
rect 13082 42469 13174 42535
rect 13082 42423 13115 42469
rect 13161 42423 13174 42469
rect 13082 42357 13174 42423
rect 13082 42311 13115 42357
rect 13161 42311 13174 42357
rect 13082 42245 13174 42311
rect 13082 42199 13115 42245
rect 13161 42199 13174 42245
rect 13082 42146 13174 42199
rect 13530 42693 13622 42746
rect 13530 42647 13543 42693
rect 13589 42647 13622 42693
rect 13530 42581 13622 42647
rect 13530 42535 13543 42581
rect 13589 42535 13622 42581
rect 13530 42469 13622 42535
rect 13530 42423 13543 42469
rect 13589 42423 13622 42469
rect 13530 42357 13622 42423
rect 13530 42311 13543 42357
rect 13589 42311 13622 42357
rect 13530 42245 13622 42311
rect 13530 42199 13543 42245
rect 13589 42199 13622 42245
rect 13530 42146 13622 42199
rect 14222 42693 14314 42746
rect 14222 42647 14255 42693
rect 14301 42647 14314 42693
rect 14222 42581 14314 42647
rect 14222 42535 14255 42581
rect 14301 42535 14314 42581
rect 14222 42469 14314 42535
rect 14222 42423 14255 42469
rect 14301 42423 14314 42469
rect 14222 42357 14314 42423
rect 14222 42311 14255 42357
rect 14301 42311 14314 42357
rect 14222 42245 14314 42311
rect 14222 42199 14255 42245
rect 14301 42199 14314 42245
rect 14222 42146 14314 42199
rect 12390 41725 12482 41778
rect 12390 41679 12403 41725
rect 12449 41679 12482 41725
rect 12390 41613 12482 41679
rect 12390 41567 12403 41613
rect 12449 41567 12482 41613
rect 12390 41501 12482 41567
rect 12390 41455 12403 41501
rect 12449 41455 12482 41501
rect 12390 41389 12482 41455
rect 12390 41343 12403 41389
rect 12449 41343 12482 41389
rect 12390 41277 12482 41343
rect 12390 41231 12403 41277
rect 12449 41231 12482 41277
rect 12390 41178 12482 41231
rect 13082 41725 13174 41778
rect 13082 41679 13115 41725
rect 13161 41679 13174 41725
rect 13082 41613 13174 41679
rect 13082 41567 13115 41613
rect 13161 41567 13174 41613
rect 13082 41501 13174 41567
rect 13082 41455 13115 41501
rect 13161 41455 13174 41501
rect 13082 41389 13174 41455
rect 13082 41343 13115 41389
rect 13161 41343 13174 41389
rect 13082 41277 13174 41343
rect 13082 41231 13115 41277
rect 13161 41231 13174 41277
rect 13082 41178 13174 41231
rect 13530 41725 13622 41778
rect 13530 41679 13543 41725
rect 13589 41679 13622 41725
rect 13530 41613 13622 41679
rect 13530 41567 13543 41613
rect 13589 41567 13622 41613
rect 13530 41501 13622 41567
rect 13530 41455 13543 41501
rect 13589 41455 13622 41501
rect 13530 41389 13622 41455
rect 13530 41343 13543 41389
rect 13589 41343 13622 41389
rect 13530 41277 13622 41343
rect 13530 41231 13543 41277
rect 13589 41231 13622 41277
rect 13530 41178 13622 41231
rect 14222 41725 14314 41778
rect 14222 41679 14255 41725
rect 14301 41679 14314 41725
rect 14222 41613 14314 41679
rect 14222 41567 14255 41613
rect 14301 41567 14314 41613
rect 14222 41501 14314 41567
rect 14222 41455 14255 41501
rect 14301 41455 14314 41501
rect 14222 41389 14314 41455
rect 14222 41343 14255 41389
rect 14301 41343 14314 41389
rect 14222 41277 14314 41343
rect 14222 41231 14255 41277
rect 14301 41231 14314 41277
rect 14222 41178 14314 41231
<< polycontact >>
rect 2681 56320 2727 56366
rect 2681 56172 2727 56218
rect 3793 56320 3839 56366
rect 3793 56172 3839 56218
rect 4181 56320 4227 56366
rect 4181 56172 4227 56218
rect 5293 56320 5339 56366
rect 5293 56172 5339 56218
rect 5681 56320 5727 56366
rect 5681 56172 5727 56218
rect 6793 56320 6839 56366
rect 6793 56172 6839 56218
rect 7181 56320 7227 56366
rect 7181 56172 7227 56218
rect 8293 56320 8339 56366
rect 8293 56172 8339 56218
rect 8681 56320 8727 56366
rect 8681 56172 8727 56218
rect 9793 56320 9839 56366
rect 9793 56172 9839 56218
rect 10181 56320 10227 56366
rect 10181 56172 10227 56218
rect 11293 56320 11339 56366
rect 11293 56172 11339 56218
rect 11681 56320 11727 56366
rect 11681 56172 11727 56218
rect 12793 56320 12839 56366
rect 12793 56172 12839 56218
rect 13181 56320 13227 56366
rect 13181 56172 13227 56218
rect 14293 56320 14339 56366
rect 14293 56172 14339 56218
rect 1403 55485 1449 55531
rect 1403 55033 1449 55079
rect 1683 55485 1729 55531
rect 1683 55033 1729 55079
rect 12403 42647 12449 42693
rect 12403 42535 12449 42581
rect 12403 42423 12449 42469
rect 12403 42311 12449 42357
rect 12403 42199 12449 42245
rect 13115 42647 13161 42693
rect 13115 42535 13161 42581
rect 13115 42423 13161 42469
rect 13115 42311 13161 42357
rect 13115 42199 13161 42245
rect 13543 42647 13589 42693
rect 13543 42535 13589 42581
rect 13543 42423 13589 42469
rect 13543 42311 13589 42357
rect 13543 42199 13589 42245
rect 14255 42647 14301 42693
rect 14255 42535 14301 42581
rect 14255 42423 14301 42469
rect 14255 42311 14301 42357
rect 14255 42199 14301 42245
rect 12403 41679 12449 41725
rect 12403 41567 12449 41613
rect 12403 41455 12449 41501
rect 12403 41343 12449 41389
rect 12403 41231 12449 41277
rect 13115 41679 13161 41725
rect 13115 41567 13161 41613
rect 13115 41455 13161 41501
rect 13115 41343 13161 41389
rect 13115 41231 13161 41277
rect 13543 41679 13589 41725
rect 13543 41567 13589 41613
rect 13543 41455 13589 41501
rect 13543 41343 13589 41389
rect 13543 41231 13589 41277
rect 14255 41679 14301 41725
rect 14255 41567 14301 41613
rect 14255 41455 14301 41501
rect 14255 41343 14301 41389
rect 14255 41231 14301 41277
<< ppolyres >>
rect 1346 55122 1506 55442
rect 1626 55122 1786 55442
<< mvpdiode >>
rect 11458 41444 11658 41457
rect 11458 41398 11471 41444
rect 11517 41398 11599 41444
rect 11645 41398 11658 41444
rect 11458 41316 11658 41398
rect 11458 41270 11471 41316
rect 11517 41270 11599 41316
rect 11645 41270 11658 41316
rect 11458 41257 11658 41270
rect 11458 40980 11658 40993
rect 11458 40934 11471 40980
rect 11517 40934 11599 40980
rect 11645 40934 11658 40980
rect 11458 40852 11658 40934
rect 11458 40806 11471 40852
rect 11517 40806 11599 40852
rect 11645 40806 11658 40852
rect 11458 40793 11658 40806
<< mvpdiodec >>
rect 11471 41398 11517 41444
rect 11599 41398 11645 41444
rect 11471 41270 11517 41316
rect 11599 41270 11645 41316
rect 11471 40934 11517 40980
rect 11599 40934 11645 40980
rect 11471 40806 11517 40852
rect 11599 40806 11645 40852
<< metal1 >>
rect 0 52180 122 57187
rect 2342 56832 14724 56843
rect 2342 56786 2353 56832
rect 14713 56786 14724 56832
rect 2342 56738 2522 56786
rect 2574 56738 2646 56786
rect 2698 56738 2770 56786
rect 2822 56738 2894 56786
rect 2946 56738 3018 56786
rect 3070 56738 3142 56786
rect 3194 56738 3266 56786
rect 3318 56738 3390 56786
rect 3442 56738 3514 56786
rect 3566 56738 3638 56786
rect 3690 56738 3762 56786
rect 3814 56738 3886 56786
rect 3938 56738 4010 56786
rect 4062 56738 4134 56786
rect 4186 56738 4258 56786
rect 4310 56738 4382 56786
rect 4434 56738 4506 56786
rect 4558 56738 4630 56786
rect 4682 56738 4754 56786
rect 4806 56738 4878 56786
rect 4930 56738 5002 56786
rect 5054 56738 5126 56786
rect 5178 56738 5250 56786
rect 5302 56738 5374 56786
rect 5426 56738 5498 56786
rect 5550 56738 5622 56786
rect 5674 56738 5746 56786
rect 5798 56738 5870 56786
rect 5922 56738 5994 56786
rect 6046 56738 6118 56786
rect 6170 56738 6242 56786
rect 6294 56738 6366 56786
rect 6418 56738 6490 56786
rect 6542 56738 6614 56786
rect 6666 56738 6738 56786
rect 6790 56738 6862 56786
rect 6914 56738 6986 56786
rect 7038 56738 7110 56786
rect 7162 56738 7234 56786
rect 7286 56738 7358 56786
rect 7410 56738 7482 56786
rect 7534 56738 7606 56786
rect 7658 56738 7730 56786
rect 7782 56738 7854 56786
rect 7906 56738 7978 56786
rect 8030 56738 8102 56786
rect 8154 56738 8226 56786
rect 8278 56738 8350 56786
rect 8402 56738 8474 56786
rect 8526 56738 8598 56786
rect 8650 56738 8722 56786
rect 8774 56738 8846 56786
rect 8898 56738 8970 56786
rect 9022 56738 9094 56786
rect 9146 56738 9218 56786
rect 9270 56738 9342 56786
rect 9394 56738 9466 56786
rect 9518 56738 9590 56786
rect 9642 56738 9714 56786
rect 9766 56738 9838 56786
rect 9890 56738 9962 56786
rect 10014 56738 10086 56786
rect 10138 56738 10210 56786
rect 10262 56738 10334 56786
rect 10386 56738 10458 56786
rect 10510 56738 10582 56786
rect 10634 56738 10706 56786
rect 10758 56738 10830 56786
rect 10882 56738 10954 56786
rect 11006 56738 11078 56786
rect 11130 56738 11202 56786
rect 11254 56738 11326 56786
rect 11378 56738 11450 56786
rect 11502 56738 11574 56786
rect 11626 56738 11698 56786
rect 11750 56738 11822 56786
rect 11874 56738 11946 56786
rect 11998 56738 12070 56786
rect 12122 56738 12194 56786
rect 12246 56738 12318 56786
rect 12370 56738 12442 56786
rect 12494 56738 12566 56786
rect 12618 56738 12690 56786
rect 12742 56738 12814 56786
rect 12866 56738 12938 56786
rect 12990 56738 13062 56786
rect 13114 56738 13186 56786
rect 13238 56738 13310 56786
rect 13362 56738 13434 56786
rect 13486 56738 13558 56786
rect 13610 56738 14724 56786
rect 2342 56668 14724 56738
rect 2342 55870 2353 56668
rect 2399 56666 14667 56668
rect 2399 56614 2522 56666
rect 2574 56614 2646 56666
rect 2698 56614 2770 56666
rect 2822 56614 2894 56666
rect 2946 56614 3018 56666
rect 3070 56614 3142 56666
rect 3194 56614 3266 56666
rect 3318 56614 3390 56666
rect 3442 56614 3514 56666
rect 3566 56614 3638 56666
rect 3690 56614 3762 56666
rect 3814 56614 3886 56666
rect 3938 56614 4010 56666
rect 4062 56614 4134 56666
rect 4186 56614 4258 56666
rect 4310 56614 4382 56666
rect 4434 56614 4506 56666
rect 4558 56614 4630 56666
rect 4682 56614 4754 56666
rect 4806 56614 4878 56666
rect 4930 56614 5002 56666
rect 5054 56614 5126 56666
rect 5178 56614 5250 56666
rect 5302 56614 5374 56666
rect 5426 56614 5498 56666
rect 5550 56614 5622 56666
rect 5674 56614 5746 56666
rect 5798 56614 5870 56666
rect 5922 56614 5994 56666
rect 6046 56614 6118 56666
rect 6170 56614 6242 56666
rect 6294 56614 6366 56666
rect 6418 56614 6490 56666
rect 6542 56614 6614 56666
rect 6666 56614 6738 56666
rect 6790 56614 6862 56666
rect 6914 56614 6986 56666
rect 7038 56614 7110 56666
rect 7162 56614 7234 56666
rect 7286 56614 7358 56666
rect 7410 56614 7482 56666
rect 7534 56614 7606 56666
rect 7658 56614 7730 56666
rect 7782 56614 7854 56666
rect 7906 56614 7978 56666
rect 8030 56614 8102 56666
rect 8154 56614 8226 56666
rect 8278 56614 8350 56666
rect 8402 56614 8474 56666
rect 8526 56614 8598 56666
rect 8650 56614 8722 56666
rect 8774 56614 8846 56666
rect 8898 56614 8970 56666
rect 9022 56614 9094 56666
rect 9146 56614 9218 56666
rect 9270 56614 9342 56666
rect 9394 56614 9466 56666
rect 9518 56614 9590 56666
rect 9642 56614 9714 56666
rect 9766 56614 9838 56666
rect 9890 56614 9962 56666
rect 10014 56614 10086 56666
rect 10138 56614 10210 56666
rect 10262 56614 10334 56666
rect 10386 56614 10458 56666
rect 10510 56614 10582 56666
rect 10634 56614 10706 56666
rect 10758 56614 10830 56666
rect 10882 56614 10954 56666
rect 11006 56614 11078 56666
rect 11130 56614 11202 56666
rect 11254 56614 11326 56666
rect 11378 56614 11450 56666
rect 11502 56614 11574 56666
rect 11626 56614 11698 56666
rect 11750 56614 11822 56666
rect 11874 56614 11946 56666
rect 11998 56614 12070 56666
rect 12122 56614 12194 56666
rect 12246 56614 12318 56666
rect 12370 56614 12442 56666
rect 12494 56614 12566 56666
rect 12618 56614 12690 56666
rect 12742 56614 12814 56666
rect 12866 56614 12938 56666
rect 12990 56614 13062 56666
rect 13114 56614 13186 56666
rect 13238 56614 13310 56666
rect 13362 56614 13434 56666
rect 13486 56614 13558 56666
rect 13610 56614 14667 56666
rect 2399 56542 14667 56614
rect 2399 56490 2522 56542
rect 2574 56490 2646 56542
rect 2698 56490 2770 56542
rect 2822 56494 2894 56542
rect 2946 56494 3018 56542
rect 3070 56494 3142 56542
rect 3194 56494 3266 56542
rect 3318 56494 3390 56542
rect 3442 56494 3514 56542
rect 3566 56494 3638 56542
rect 3690 56494 3762 56542
rect 3723 56490 3762 56494
rect 3814 56490 3886 56542
rect 3938 56490 4010 56542
rect 4062 56490 4134 56542
rect 4186 56490 4258 56542
rect 4310 56494 4382 56542
rect 4434 56494 4506 56542
rect 4558 56494 4630 56542
rect 4682 56494 4754 56542
rect 4806 56494 4878 56542
rect 4930 56494 5002 56542
rect 5054 56494 5126 56542
rect 5178 56494 5250 56542
rect 5223 56490 5250 56494
rect 5302 56490 5374 56542
rect 5426 56490 5498 56542
rect 5550 56490 5622 56542
rect 5674 56490 5746 56542
rect 5798 56494 5870 56542
rect 5922 56494 5994 56542
rect 6046 56494 6118 56542
rect 6170 56494 6242 56542
rect 6294 56494 6366 56542
rect 6418 56494 6490 56542
rect 6542 56494 6614 56542
rect 6666 56494 6738 56542
rect 6723 56490 6738 56494
rect 6790 56490 6862 56542
rect 6914 56490 6986 56542
rect 7038 56490 7110 56542
rect 7162 56490 7234 56542
rect 7286 56494 7358 56542
rect 7410 56494 7482 56542
rect 7534 56494 7606 56542
rect 7658 56494 7730 56542
rect 7782 56494 7854 56542
rect 7906 56494 7978 56542
rect 8030 56494 8102 56542
rect 8154 56494 8226 56542
rect 7286 56490 7297 56494
rect 8223 56490 8226 56494
rect 8278 56490 8350 56542
rect 8402 56490 8474 56542
rect 8526 56490 8598 56542
rect 8650 56490 8722 56542
rect 8774 56494 8846 56542
rect 8898 56494 8970 56542
rect 9022 56494 9094 56542
rect 9146 56494 9218 56542
rect 9270 56494 9342 56542
rect 9394 56494 9466 56542
rect 9518 56494 9590 56542
rect 9642 56494 9714 56542
rect 8774 56490 8797 56494
rect 9766 56490 9838 56542
rect 9890 56490 9962 56542
rect 10014 56490 10086 56542
rect 10138 56490 10210 56542
rect 10262 56494 10334 56542
rect 10386 56494 10458 56542
rect 10510 56494 10582 56542
rect 10634 56494 10706 56542
rect 10758 56494 10830 56542
rect 10882 56494 10954 56542
rect 11006 56494 11078 56542
rect 11130 56494 11202 56542
rect 10262 56490 10297 56494
rect 11254 56490 11326 56542
rect 11378 56490 11450 56542
rect 11502 56490 11574 56542
rect 11626 56490 11698 56542
rect 11750 56494 11822 56542
rect 11874 56494 11946 56542
rect 11998 56494 12070 56542
rect 12122 56494 12194 56542
rect 12246 56494 12318 56542
rect 12370 56494 12442 56542
rect 12494 56494 12566 56542
rect 12618 56494 12690 56542
rect 11750 56490 11797 56494
rect 12742 56490 12814 56542
rect 12866 56490 12938 56542
rect 12990 56490 13062 56542
rect 13114 56490 13186 56542
rect 13238 56494 13310 56542
rect 13362 56494 13434 56542
rect 13486 56494 13558 56542
rect 13610 56494 14667 56542
rect 13238 56490 13297 56494
rect 2399 56448 2797 56490
rect 3723 56448 4297 56490
rect 5223 56448 5797 56490
rect 6723 56448 7297 56490
rect 8223 56448 8797 56490
rect 9723 56448 10297 56490
rect 11223 56448 11797 56490
rect 12723 56448 13297 56490
rect 14223 56448 14667 56494
rect 2399 56437 14667 56448
rect 2399 56101 2610 56437
rect 2670 56366 3850 56377
rect 2670 56320 2681 56366
rect 2727 56345 3793 56366
rect 2670 56218 2682 56320
rect 2670 56172 2681 56218
rect 2838 56189 3682 56345
rect 3839 56320 3850 56366
rect 3838 56218 3850 56320
rect 2727 56172 3793 56189
rect 3839 56172 3850 56218
rect 2670 56161 3850 56172
rect 3910 56101 4110 56437
rect 4170 56366 5350 56377
rect 4170 56320 4181 56366
rect 4227 56345 5293 56366
rect 4170 56218 4182 56320
rect 4170 56172 4181 56218
rect 4338 56189 5182 56345
rect 5339 56320 5350 56366
rect 5338 56218 5350 56320
rect 4227 56172 5293 56189
rect 5339 56172 5350 56218
rect 4170 56161 5350 56172
rect 5410 56101 5610 56437
rect 5670 56366 6850 56377
rect 5670 56320 5681 56366
rect 5727 56345 6793 56366
rect 5670 56218 5682 56320
rect 5670 56172 5681 56218
rect 5838 56189 6682 56345
rect 6839 56320 6850 56366
rect 6838 56218 6850 56320
rect 5727 56172 6793 56189
rect 6839 56172 6850 56218
rect 5670 56161 6850 56172
rect 6910 56101 7110 56437
rect 7170 56366 8350 56377
rect 7170 56320 7181 56366
rect 7227 56345 8293 56366
rect 7170 56218 7182 56320
rect 7170 56172 7181 56218
rect 7338 56189 8182 56345
rect 8339 56320 8350 56366
rect 8338 56218 8350 56320
rect 7227 56172 8293 56189
rect 8339 56172 8350 56218
rect 7170 56161 8350 56172
rect 8410 56101 8610 56437
rect 8670 56366 9850 56377
rect 8670 56320 8681 56366
rect 8727 56345 9793 56366
rect 8670 56218 8682 56320
rect 8670 56172 8681 56218
rect 8838 56189 9682 56345
rect 9839 56320 9850 56366
rect 9838 56218 9850 56320
rect 8727 56172 9793 56189
rect 9839 56172 9850 56218
rect 8670 56161 9850 56172
rect 9910 56101 10110 56437
rect 10170 56366 11350 56377
rect 10170 56320 10181 56366
rect 10227 56345 11293 56366
rect 10170 56218 10182 56320
rect 10170 56172 10181 56218
rect 10338 56189 11182 56345
rect 11339 56320 11350 56366
rect 11338 56218 11350 56320
rect 10227 56172 11293 56189
rect 11339 56172 11350 56218
rect 10170 56161 11350 56172
rect 11410 56101 11610 56437
rect 11670 56366 12850 56377
rect 11670 56320 11681 56366
rect 11727 56345 12793 56366
rect 11670 56218 11682 56320
rect 11670 56172 11681 56218
rect 11838 56189 12682 56345
rect 12839 56320 12850 56366
rect 12838 56218 12850 56320
rect 11727 56172 12793 56189
rect 12839 56172 12850 56218
rect 11670 56161 12850 56172
rect 12910 56101 13110 56437
rect 13170 56366 14560 56377
rect 13170 56320 13181 56366
rect 13227 56345 14293 56366
rect 13338 56320 14293 56345
rect 14339 56345 14560 56366
rect 14339 56320 14392 56345
rect 13170 56218 13182 56320
rect 13338 56218 14392 56320
rect 13170 56172 13181 56218
rect 13338 56189 14293 56218
rect 13227 56172 14293 56189
rect 14339 56189 14392 56218
rect 14548 56189 14560 56345
rect 14339 56172 14560 56189
rect 13170 56161 14560 56172
rect 14656 56101 14667 56437
rect 2399 56090 14667 56101
rect 2399 56048 2797 56090
rect 3723 56048 4297 56090
rect 5223 56048 5797 56090
rect 6723 56048 7297 56090
rect 8223 56048 8797 56090
rect 9723 56048 10297 56090
rect 11223 56048 11797 56090
rect 12723 56048 13297 56090
rect 2399 55996 2522 56048
rect 2574 55996 2646 56048
rect 2698 55996 2770 56048
rect 3723 56044 3762 56048
rect 2822 55996 2894 56044
rect 2946 55996 3018 56044
rect 3070 55996 3142 56044
rect 3194 55996 3266 56044
rect 3318 55996 3390 56044
rect 3442 55996 3514 56044
rect 3566 55996 3638 56044
rect 3690 55996 3762 56044
rect 3814 55996 3886 56048
rect 3938 55996 4010 56048
rect 4062 55996 4134 56048
rect 4186 55996 4258 56048
rect 5223 56044 5250 56048
rect 4310 55996 4382 56044
rect 4434 55996 4506 56044
rect 4558 55996 4630 56044
rect 4682 55996 4754 56044
rect 4806 55996 4878 56044
rect 4930 55996 5002 56044
rect 5054 55996 5126 56044
rect 5178 55996 5250 56044
rect 5302 55996 5374 56048
rect 5426 55996 5498 56048
rect 5550 55996 5622 56048
rect 5674 55996 5746 56048
rect 6723 56044 6738 56048
rect 5798 55996 5870 56044
rect 5922 55996 5994 56044
rect 6046 55996 6118 56044
rect 6170 55996 6242 56044
rect 6294 55996 6366 56044
rect 6418 55996 6490 56044
rect 6542 55996 6614 56044
rect 6666 55996 6738 56044
rect 6790 55996 6862 56048
rect 6914 55996 6986 56048
rect 7038 55996 7110 56048
rect 7162 55996 7234 56048
rect 7286 56044 7297 56048
rect 8223 56044 8226 56048
rect 7286 55996 7358 56044
rect 7410 55996 7482 56044
rect 7534 55996 7606 56044
rect 7658 55996 7730 56044
rect 7782 55996 7854 56044
rect 7906 55996 7978 56044
rect 8030 55996 8102 56044
rect 8154 55996 8226 56044
rect 8278 55996 8350 56048
rect 8402 55996 8474 56048
rect 8526 55996 8598 56048
rect 8650 55996 8722 56048
rect 8774 56044 8797 56048
rect 8774 55996 8846 56044
rect 8898 55996 8970 56044
rect 9022 55996 9094 56044
rect 9146 55996 9218 56044
rect 9270 55996 9342 56044
rect 9394 55996 9466 56044
rect 9518 55996 9590 56044
rect 9642 55996 9714 56044
rect 9766 55996 9838 56048
rect 9890 55996 9962 56048
rect 10014 55996 10086 56048
rect 10138 55996 10210 56048
rect 10262 56044 10297 56048
rect 10262 55996 10334 56044
rect 10386 55996 10458 56044
rect 10510 55996 10582 56044
rect 10634 55996 10706 56044
rect 10758 55996 10830 56044
rect 10882 55996 10954 56044
rect 11006 55996 11078 56044
rect 11130 55996 11202 56044
rect 11254 55996 11326 56048
rect 11378 55996 11450 56048
rect 11502 55996 11574 56048
rect 11626 55996 11698 56048
rect 11750 56044 11797 56048
rect 11750 55996 11822 56044
rect 11874 55996 11946 56044
rect 11998 55996 12070 56044
rect 12122 55996 12194 56044
rect 12246 55996 12318 56044
rect 12370 55996 12442 56044
rect 12494 55996 12566 56044
rect 12618 55996 12690 56044
rect 12742 55996 12814 56048
rect 12866 55996 12938 56048
rect 12990 55996 13062 56048
rect 13114 55996 13186 56048
rect 13238 56044 13297 56048
rect 14223 56044 14667 56090
rect 13238 55996 13310 56044
rect 13362 55996 13434 56044
rect 13486 55996 13558 56044
rect 13610 55996 14667 56044
rect 2399 55924 14667 55996
rect 2399 55872 2522 55924
rect 2574 55872 2646 55924
rect 2698 55872 2770 55924
rect 2822 55872 2894 55924
rect 2946 55872 3018 55924
rect 3070 55872 3142 55924
rect 3194 55872 3266 55924
rect 3318 55872 3390 55924
rect 3442 55872 3514 55924
rect 3566 55872 3638 55924
rect 3690 55872 3762 55924
rect 3814 55872 3886 55924
rect 3938 55872 4010 55924
rect 4062 55872 4134 55924
rect 4186 55872 4258 55924
rect 4310 55872 4382 55924
rect 4434 55872 4506 55924
rect 4558 55872 4630 55924
rect 4682 55872 4754 55924
rect 4806 55872 4878 55924
rect 4930 55872 5002 55924
rect 5054 55872 5126 55924
rect 5178 55872 5250 55924
rect 5302 55872 5374 55924
rect 5426 55872 5498 55924
rect 5550 55872 5622 55924
rect 5674 55872 5746 55924
rect 5798 55872 5870 55924
rect 5922 55872 5994 55924
rect 6046 55872 6118 55924
rect 6170 55872 6242 55924
rect 6294 55872 6366 55924
rect 6418 55872 6490 55924
rect 6542 55872 6614 55924
rect 6666 55872 6738 55924
rect 6790 55872 6862 55924
rect 6914 55872 6986 55924
rect 7038 55872 7110 55924
rect 7162 55872 7234 55924
rect 7286 55872 7358 55924
rect 7410 55872 7482 55924
rect 7534 55872 7606 55924
rect 7658 55872 7730 55924
rect 7782 55872 7854 55924
rect 7906 55872 7978 55924
rect 8030 55872 8102 55924
rect 8154 55872 8226 55924
rect 8278 55872 8350 55924
rect 8402 55872 8474 55924
rect 8526 55872 8598 55924
rect 8650 55872 8722 55924
rect 8774 55872 8846 55924
rect 8898 55872 8970 55924
rect 9022 55872 9094 55924
rect 9146 55872 9218 55924
rect 9270 55872 9342 55924
rect 9394 55872 9466 55924
rect 9518 55872 9590 55924
rect 9642 55872 9714 55924
rect 9766 55872 9838 55924
rect 9890 55872 9962 55924
rect 10014 55872 10086 55924
rect 10138 55872 10210 55924
rect 10262 55872 10334 55924
rect 10386 55872 10458 55924
rect 10510 55872 10582 55924
rect 10634 55872 10706 55924
rect 10758 55872 10830 55924
rect 10882 55872 10954 55924
rect 11006 55872 11078 55924
rect 11130 55872 11202 55924
rect 11254 55872 11326 55924
rect 11378 55872 11450 55924
rect 11502 55872 11574 55924
rect 11626 55872 11698 55924
rect 11750 55872 11822 55924
rect 11874 55872 11946 55924
rect 11998 55872 12070 55924
rect 12122 55872 12194 55924
rect 12246 55872 12318 55924
rect 12370 55872 12442 55924
rect 12494 55872 12566 55924
rect 12618 55872 12690 55924
rect 12742 55872 12814 55924
rect 12866 55872 12938 55924
rect 12990 55872 13062 55924
rect 13114 55872 13186 55924
rect 13238 55872 13310 55924
rect 13362 55872 13434 55924
rect 13486 55872 13558 55924
rect 13610 55872 14667 55924
rect 2399 55870 14667 55872
rect 14713 55870 14724 56668
rect 1049 55822 2083 55833
rect 184 54725 921 54799
rect 1049 54742 1060 55822
rect 1106 55776 1214 55822
rect 1918 55776 2026 55822
rect 1106 55765 2026 55776
rect 1106 55090 1117 55765
rect 1348 55531 1530 55542
rect 1348 55485 1403 55531
rect 1449 55530 1530 55531
rect 1449 55485 1466 55530
rect 1348 55474 1466 55485
rect 1454 55374 1466 55474
rect 1518 55374 1530 55530
rect 1454 55362 1530 55374
rect 1596 55531 1784 55542
rect 1596 55530 1683 55531
rect 1596 55374 1608 55530
rect 1660 55485 1683 55530
rect 1729 55485 1784 55531
rect 1660 55474 1784 55485
rect 1660 55374 1672 55474
rect 1596 55362 1672 55374
rect 2015 55090 2026 55765
rect 1106 55079 2026 55090
rect 1106 55033 1403 55079
rect 1449 55033 1683 55079
rect 1729 55033 2026 55079
rect 1106 55022 2026 55033
rect 1106 54742 1117 55022
rect 1049 54731 1117 54742
rect 1203 54788 1929 54799
rect 1203 54742 1214 54788
rect 1918 54742 1929 54788
rect 1203 54731 1929 54742
rect 2015 54742 2026 55022
rect 2072 54742 2083 55822
rect 2342 55800 14724 55870
rect 2342 55752 2522 55800
rect 2574 55752 2646 55800
rect 2698 55752 2770 55800
rect 2822 55752 2894 55800
rect 2946 55752 3018 55800
rect 3070 55752 3142 55800
rect 3194 55752 3266 55800
rect 3318 55752 3390 55800
rect 3442 55752 3514 55800
rect 3566 55752 3638 55800
rect 3690 55752 3762 55800
rect 3814 55752 3886 55800
rect 3938 55752 4010 55800
rect 4062 55752 4134 55800
rect 4186 55752 4258 55800
rect 4310 55752 4382 55800
rect 4434 55752 4506 55800
rect 4558 55752 4630 55800
rect 4682 55752 4754 55800
rect 4806 55752 4878 55800
rect 4930 55752 5002 55800
rect 5054 55752 5126 55800
rect 5178 55752 5250 55800
rect 5302 55752 5374 55800
rect 5426 55752 5498 55800
rect 5550 55752 5622 55800
rect 5674 55752 5746 55800
rect 5798 55752 5870 55800
rect 5922 55752 5994 55800
rect 6046 55752 6118 55800
rect 6170 55752 6242 55800
rect 6294 55752 6366 55800
rect 6418 55752 6490 55800
rect 6542 55752 6614 55800
rect 6666 55752 6738 55800
rect 6790 55752 6862 55800
rect 6914 55752 6986 55800
rect 7038 55752 7110 55800
rect 7162 55752 7234 55800
rect 7286 55752 7358 55800
rect 7410 55752 7482 55800
rect 7534 55752 7606 55800
rect 7658 55752 7730 55800
rect 7782 55752 7854 55800
rect 7906 55752 7978 55800
rect 8030 55752 8102 55800
rect 8154 55752 8226 55800
rect 8278 55752 8350 55800
rect 8402 55752 8474 55800
rect 8526 55752 8598 55800
rect 8650 55752 8722 55800
rect 8774 55752 8846 55800
rect 8898 55752 8970 55800
rect 9022 55752 9094 55800
rect 9146 55752 9218 55800
rect 9270 55752 9342 55800
rect 9394 55752 9466 55800
rect 9518 55752 9590 55800
rect 9642 55752 9714 55800
rect 9766 55752 9838 55800
rect 9890 55752 9962 55800
rect 10014 55752 10086 55800
rect 10138 55752 10210 55800
rect 10262 55752 10334 55800
rect 10386 55752 10458 55800
rect 10510 55752 10582 55800
rect 10634 55752 10706 55800
rect 10758 55752 10830 55800
rect 10882 55752 10954 55800
rect 11006 55752 11078 55800
rect 11130 55752 11202 55800
rect 11254 55752 11326 55800
rect 11378 55752 11450 55800
rect 11502 55752 11574 55800
rect 11626 55752 11698 55800
rect 11750 55752 11822 55800
rect 11874 55752 11946 55800
rect 11998 55752 12070 55800
rect 12122 55752 12194 55800
rect 12246 55752 12318 55800
rect 12370 55752 12442 55800
rect 12494 55752 12566 55800
rect 12618 55752 12690 55800
rect 12742 55752 12814 55800
rect 12866 55752 12938 55800
rect 12990 55752 13062 55800
rect 13114 55752 13186 55800
rect 13238 55752 13310 55800
rect 13362 55752 13434 55800
rect 13486 55752 13558 55800
rect 13610 55752 14724 55800
rect 2342 55706 2353 55752
rect 14713 55706 14724 55752
rect 2342 55695 14724 55706
rect 2015 54731 2083 54742
rect 3470 55459 3546 55471
rect 184 54673 234 54725
rect 286 54673 358 54725
rect 410 54673 482 54725
rect 534 54673 921 54725
rect 184 54601 921 54673
rect 184 54549 234 54601
rect 286 54549 358 54601
rect 410 54549 482 54601
rect 534 54549 921 54601
rect 184 54477 921 54549
rect 184 54425 234 54477
rect 286 54425 358 54477
rect 410 54425 482 54477
rect 534 54425 921 54477
rect 3470 54471 3482 55459
rect 3534 54471 3546 55459
rect 3470 54459 3546 54471
rect 3693 55459 3769 55471
rect 3693 54471 3705 55459
rect 3757 54471 3769 55459
rect 3693 54459 3769 54471
rect 4162 55459 4238 55471
rect 4162 54471 4174 55459
rect 4226 54471 4238 55459
rect 8030 55459 8106 55471
rect 4758 55404 4834 55416
rect 4758 54624 4770 55404
rect 4822 54624 4834 55404
rect 4758 54612 4834 54624
rect 4938 55404 5014 55416
rect 4938 54624 4950 55404
rect 5002 54624 5014 55404
rect 4938 54612 5014 54624
rect 5426 55404 5502 55416
rect 5426 54624 5438 55404
rect 5490 54624 5502 55404
rect 5426 54612 5502 54624
rect 5914 55404 5990 55416
rect 5914 54624 5926 55404
rect 5978 54624 5990 55404
rect 6278 55404 6354 55416
rect 5914 54612 5990 54624
rect 6096 55359 6172 55403
rect 4162 54459 4238 54471
rect 6096 54475 6108 55359
rect 6160 54475 6172 55359
rect 6278 54624 6290 55404
rect 6342 54624 6354 55404
rect 6278 54612 6354 54624
rect 6766 55404 6842 55416
rect 6766 54624 6778 55404
rect 6830 54624 6842 55404
rect 6766 54612 6842 54624
rect 7254 55404 7330 55416
rect 7254 54624 7266 55404
rect 7318 54624 7330 55404
rect 7254 54612 7330 54624
rect 7434 55404 7510 55416
rect 7434 54624 7446 55404
rect 7498 54624 7510 55404
rect 7434 54612 7510 54624
rect 6096 54463 6172 54475
rect 8030 54471 8042 55459
rect 8094 54471 8106 55459
rect 8030 54459 8106 54471
rect 8499 55459 8575 55471
rect 8499 54471 8511 55459
rect 8563 54471 8575 55459
rect 8499 54459 8575 54471
rect 8714 55459 8790 55471
rect 8714 54471 8726 55459
rect 8778 54471 8790 55459
rect 8714 54459 8790 54471
rect 8937 55459 9013 55471
rect 8937 54471 8949 55459
rect 9001 54471 9013 55459
rect 8937 54459 9013 54471
rect 9406 55459 9482 55471
rect 9406 54471 9418 55459
rect 9470 54471 9482 55459
rect 13274 55459 13350 55471
rect 10002 55404 10078 55416
rect 10002 54624 10014 55404
rect 10066 54624 10078 55404
rect 10002 54612 10078 54624
rect 10182 55404 10258 55416
rect 10182 54624 10194 55404
rect 10246 54624 10258 55404
rect 10182 54612 10258 54624
rect 10670 55404 10746 55416
rect 10670 54624 10682 55404
rect 10734 54624 10746 55404
rect 10670 54612 10746 54624
rect 11158 55404 11234 55416
rect 11158 54624 11170 55404
rect 11222 54624 11234 55404
rect 11522 55404 11598 55416
rect 11158 54612 11234 54624
rect 11340 55359 11416 55403
rect 9406 54459 9482 54471
rect 11340 54475 11352 55359
rect 11404 54475 11416 55359
rect 11522 54624 11534 55404
rect 11586 54624 11598 55404
rect 11522 54612 11598 54624
rect 12010 55404 12086 55416
rect 12010 54624 12022 55404
rect 12074 54624 12086 55404
rect 12010 54612 12086 54624
rect 12498 55404 12574 55416
rect 12498 54624 12510 55404
rect 12562 54624 12574 55404
rect 12498 54612 12574 54624
rect 12678 55404 12754 55416
rect 12678 54624 12690 55404
rect 12742 54624 12754 55404
rect 12678 54612 12754 54624
rect 11340 54463 11416 54475
rect 13274 54471 13286 55459
rect 13338 54471 13350 55459
rect 13274 54459 13350 54471
rect 184 54354 921 54425
rect 3470 54001 3546 54013
rect 184 53825 921 53890
rect 184 53773 234 53825
rect 286 53773 358 53825
rect 410 53773 482 53825
rect 534 53773 921 53825
rect 184 53701 921 53773
rect 184 53649 234 53701
rect 286 53649 358 53701
rect 410 53649 482 53701
rect 534 53649 921 53701
rect 184 53577 921 53649
rect 184 53525 234 53577
rect 286 53525 358 53577
rect 410 53525 482 53577
rect 534 53525 921 53577
rect 184 53454 921 53525
rect 3470 53013 3482 54001
rect 3534 53013 3546 54001
rect 8718 54001 8794 54013
rect 6096 53897 6172 53909
rect 3470 53001 3546 53013
rect 4162 53793 4238 53805
rect 4162 53013 4174 53793
rect 4226 53013 4238 53793
rect 4758 53632 4834 53644
rect 4758 53060 4770 53632
rect 4822 53060 4834 53632
rect 4758 53048 4834 53060
rect 4938 53632 5014 53644
rect 4938 53060 4950 53632
rect 5002 53060 5014 53632
rect 4938 53048 5014 53060
rect 5426 53632 5502 53644
rect 5426 53060 5438 53632
rect 5490 53060 5502 53632
rect 5426 53048 5502 53060
rect 5914 53632 5990 53644
rect 5914 53060 5926 53632
rect 5978 53060 5990 53632
rect 5914 53048 5990 53060
rect 4162 53001 4238 53013
rect 6096 53013 6108 53897
rect 6160 53013 6172 53897
rect 8030 53793 8106 53805
rect 6278 53632 6354 53644
rect 6278 53060 6290 53632
rect 6342 53060 6354 53632
rect 6278 53048 6354 53060
rect 6766 53632 6842 53644
rect 6766 53060 6778 53632
rect 6830 53060 6842 53632
rect 6766 53048 6842 53060
rect 7254 53632 7330 53644
rect 7254 53060 7266 53632
rect 7318 53060 7330 53632
rect 7254 53048 7330 53060
rect 7434 53632 7510 53644
rect 7434 53060 7446 53632
rect 7498 53060 7510 53632
rect 7434 53048 7510 53060
rect 6096 53001 6172 53013
rect 8030 53013 8042 53793
rect 8094 53013 8106 53793
rect 8030 53001 8106 53013
rect 8718 53013 8730 54001
rect 8782 53013 8794 54001
rect 11340 53897 11416 53909
rect 10002 53632 10078 53644
rect 10002 53060 10014 53632
rect 10066 53060 10078 53632
rect 10002 53048 10078 53060
rect 10182 53632 10258 53644
rect 10182 53060 10194 53632
rect 10246 53060 10258 53632
rect 10182 53048 10258 53060
rect 10670 53632 10746 53644
rect 10670 53060 10682 53632
rect 10734 53060 10746 53632
rect 10670 53048 10746 53060
rect 11158 53632 11234 53644
rect 11158 53060 11170 53632
rect 11222 53060 11234 53632
rect 11158 53048 11234 53060
rect 8718 53001 8794 53013
rect 11340 53013 11352 53897
rect 11404 53013 11416 53897
rect 13274 53793 13350 53805
rect 11522 53632 11598 53644
rect 11522 53060 11534 53632
rect 11586 53060 11598 53632
rect 11522 53048 11598 53060
rect 12010 53632 12086 53644
rect 12010 53060 12022 53632
rect 12074 53060 12086 53632
rect 12010 53048 12086 53060
rect 12498 53632 12574 53644
rect 12498 53060 12510 53632
rect 12562 53060 12574 53632
rect 12498 53048 12574 53060
rect 12678 53632 12754 53644
rect 12678 53060 12690 53632
rect 12742 53060 12754 53632
rect 12678 53048 12754 53060
rect 11340 53001 11416 53013
rect 13274 53013 13286 53793
rect 13338 53013 13350 53793
rect 13274 53001 13350 53013
rect 704 52637 3895 52649
rect 704 52585 722 52637
rect 1086 52585 3378 52637
rect 3534 52585 3727 52637
rect 3883 52585 3895 52637
rect 704 52573 3895 52585
rect 6438 52309 6930 52321
rect 6438 52257 6450 52309
rect 6918 52257 6930 52309
rect 6438 52245 6930 52257
rect 7254 52309 7434 52321
rect 7254 52257 7266 52309
rect 7422 52257 7434 52309
rect 7254 52245 7434 52257
rect 0 50880 58 52180
rect 110 50880 122 52180
rect 0 37780 122 50880
rect 14942 52180 15064 57187
rect 14942 50880 14954 52180
rect 15006 50880 15064 52180
rect 2528 49899 6140 49911
rect 2528 49847 2540 49899
rect 6128 49847 6140 49899
rect 2528 49835 6140 49847
rect 7720 49899 8108 49911
rect 7720 49847 7732 49899
rect 8096 49847 8108 49899
rect 7720 49835 8108 49847
rect 8422 49899 8810 49911
rect 8422 49847 8434 49899
rect 8798 49847 8810 49899
rect 8422 49835 8810 49847
rect 4632 49054 4956 49066
rect 3904 48916 4366 49030
rect 3904 48864 3990 48916
rect 4042 48864 4114 48916
rect 4166 48864 4238 48916
rect 4290 48864 4366 48916
rect 3904 48792 4366 48864
rect 3904 48740 3990 48792
rect 4042 48740 4114 48792
rect 4166 48740 4238 48792
rect 4290 48740 4366 48792
rect 3904 48668 4366 48740
rect 3904 48616 3990 48668
rect 4042 48616 4114 48668
rect 4166 48616 4238 48668
rect 4290 48616 4366 48668
rect 3904 48544 4366 48616
rect 3904 48492 3990 48544
rect 4042 48492 4114 48544
rect 4166 48492 4238 48544
rect 4290 48492 4366 48544
rect 3904 48420 4366 48492
rect 3904 48368 3990 48420
rect 4042 48368 4114 48420
rect 4166 48368 4238 48420
rect 4290 48368 4366 48420
rect 3904 48296 4366 48368
rect 3904 48244 3990 48296
rect 4042 48244 4114 48296
rect 4166 48244 4238 48296
rect 4290 48244 4366 48296
rect 3904 48172 4366 48244
rect 3904 48120 3990 48172
rect 4042 48120 4114 48172
rect 4166 48120 4238 48172
rect 4290 48120 4366 48172
rect 3904 48048 4366 48120
rect 3904 47996 3990 48048
rect 4042 47996 4114 48048
rect 4166 47996 4238 48048
rect 4290 47996 4366 48048
rect 3904 47924 4366 47996
rect 3904 47872 3990 47924
rect 4042 47872 4114 47924
rect 4166 47872 4238 47924
rect 4290 47872 4366 47924
rect 3904 47800 4366 47872
rect 3904 47748 3990 47800
rect 4042 47748 4114 47800
rect 4166 47748 4238 47800
rect 4290 47748 4366 47800
rect 3608 47418 3684 47430
rect 3608 46326 3620 47418
rect 3672 46326 3684 47418
rect 3608 46314 3684 46326
rect 3185 46134 3365 46150
rect 3185 45666 3197 46134
rect 3353 45666 3365 46134
rect 3185 45654 3365 45666
rect 3904 45339 4366 47748
rect 4632 49002 4644 49054
rect 4696 49002 4768 49054
rect 4820 49002 4892 49054
rect 4944 49002 4956 49054
rect 4632 48930 4956 49002
rect 4632 48878 4644 48930
rect 4696 48878 4768 48930
rect 4820 48878 4892 48930
rect 4944 48878 4956 48930
rect 4632 48806 4956 48878
rect 4632 48754 4644 48806
rect 4696 48754 4768 48806
rect 4820 48754 4892 48806
rect 4944 48754 4956 48806
rect 5519 49028 5907 49040
rect 5519 48768 5531 49028
rect 5895 48768 5907 49028
rect 5519 48756 5907 48768
rect 7720 49028 8108 49040
rect 7720 48768 7732 49028
rect 8096 48768 8108 49028
rect 7720 48756 8108 48768
rect 8422 49028 8810 49040
rect 8422 48768 8434 49028
rect 8798 48768 8810 49028
rect 8422 48756 8810 48768
rect 10782 48990 10858 49002
rect 4632 48682 4956 48754
rect 4632 48630 4644 48682
rect 4696 48630 4768 48682
rect 4820 48630 4892 48682
rect 4944 48630 4956 48682
rect 4632 48558 4956 48630
rect 4632 48506 4644 48558
rect 4696 48506 4768 48558
rect 4820 48506 4892 48558
rect 4944 48506 4956 48558
rect 4632 48434 4956 48506
rect 4632 48382 4644 48434
rect 4696 48382 4768 48434
rect 4820 48382 4892 48434
rect 4944 48382 4956 48434
rect 4632 48310 4956 48382
rect 4632 48258 4644 48310
rect 4696 48258 4768 48310
rect 4820 48258 4892 48310
rect 4944 48258 4956 48310
rect 4632 48186 4956 48258
rect 4632 48134 4644 48186
rect 4696 48134 4768 48186
rect 4820 48134 4892 48186
rect 4944 48134 4956 48186
rect 4632 48062 4956 48134
rect 4632 48010 4644 48062
rect 4696 48010 4768 48062
rect 4820 48010 4892 48062
rect 4944 48010 4956 48062
rect 4632 47938 4956 48010
rect 10782 48002 10794 48990
rect 10846 48002 10858 48990
rect 10782 47990 10858 48002
rect 4632 47886 4644 47938
rect 4696 47886 4768 47938
rect 4820 47886 4892 47938
rect 4944 47886 4956 47938
rect 4632 47814 4956 47886
rect 4632 47762 4644 47814
rect 4696 47762 4768 47814
rect 4820 47762 4892 47814
rect 4944 47762 4956 47814
rect 4632 47690 4956 47762
rect 4632 47638 4644 47690
rect 4696 47638 4768 47690
rect 4820 47638 4892 47690
rect 4944 47638 4956 47690
rect 4632 47566 4956 47638
rect 4632 47514 4644 47566
rect 4696 47514 4768 47566
rect 4820 47514 4892 47566
rect 4944 47514 4956 47566
rect 4632 47502 4956 47514
rect 11567 47608 11720 47620
rect 11567 47452 11608 47608
rect 11660 47452 11720 47608
rect 11001 47404 11077 47416
rect 11001 46624 11013 47404
rect 11065 46624 11077 47404
rect 11001 46612 11077 46624
rect 11567 46092 11720 47452
rect 12002 46097 13567 46554
rect 3904 45287 3981 45339
rect 4033 45287 4105 45339
rect 4157 45287 4229 45339
rect 4281 45287 4366 45339
rect 3904 45215 4366 45287
rect 3904 45163 3981 45215
rect 4033 45163 4105 45215
rect 4157 45163 4229 45215
rect 4281 45163 4366 45215
rect 3904 45091 4366 45163
rect 3904 45039 3981 45091
rect 4033 45039 4105 45091
rect 4157 45039 4229 45091
rect 4281 45039 4366 45091
rect 3904 44967 4366 45039
rect 3904 44915 3981 44967
rect 4033 44915 4105 44967
rect 4157 44915 4229 44967
rect 4281 44915 4366 44967
rect 3904 44843 4366 44915
rect 3904 44791 3981 44843
rect 4033 44791 4105 44843
rect 4157 44791 4229 44843
rect 4281 44791 4366 44843
rect 3904 44719 4366 44791
rect 3904 44667 3981 44719
rect 4033 44667 4105 44719
rect 4157 44667 4229 44719
rect 4281 44667 4366 44719
rect 3904 44595 4366 44667
rect 3904 44543 3981 44595
rect 4033 44543 4105 44595
rect 4157 44543 4229 44595
rect 4281 44543 4366 44595
rect 3904 44430 4366 44543
rect 3608 44180 3684 44192
rect 3608 42880 3620 44180
rect 3672 42880 3684 44180
rect 12425 43683 12605 43695
rect 12425 43631 12437 43683
rect 12593 43631 12605 43683
rect 12425 43619 12605 43631
rect 3608 42868 3684 42880
rect 10470 43258 11847 43269
rect 10470 43212 10764 43258
rect 10810 43212 10878 43258
rect 10924 43212 10992 43258
rect 11038 43212 11106 43258
rect 11152 43212 11220 43258
rect 11266 43212 11334 43258
rect 11380 43212 11448 43258
rect 11494 43212 11562 43258
rect 11608 43212 11676 43258
rect 11722 43212 11790 43258
rect 11836 43218 11847 43258
rect 11836 43212 14745 43218
rect 10470 43207 14745 43212
rect 10470 43144 12075 43207
rect 10470 43098 10764 43144
rect 10810 43098 10878 43144
rect 10924 43098 10992 43144
rect 11038 43098 11106 43144
rect 11152 43098 11220 43144
rect 11266 43098 11334 43144
rect 11380 43098 11448 43144
rect 11494 43098 11562 43144
rect 11608 43098 11676 43144
rect 11722 43098 11790 43144
rect 11836 43098 12075 43144
rect 10470 43030 12075 43098
rect 10470 42984 10764 43030
rect 10810 42984 10878 43030
rect 10924 42984 10992 43030
rect 11038 42984 11106 43030
rect 11152 42984 11220 43030
rect 11266 42984 11334 43030
rect 11380 42984 11448 43030
rect 11494 42984 11562 43030
rect 11608 42984 11676 43030
rect 11722 42984 11790 43030
rect 11836 42984 12075 43030
rect 10470 42916 12075 42984
rect 10470 42870 10764 42916
rect 10810 42870 10878 42916
rect 10924 42870 10992 42916
rect 11038 42870 11106 42916
rect 11152 42870 11220 42916
rect 11266 42870 11334 42916
rect 11380 42870 11448 42916
rect 11494 42870 11562 42916
rect 11608 42870 11676 42916
rect 11722 42870 11790 42916
rect 11836 42870 12075 42916
rect 10470 42802 12075 42870
rect 10470 42773 10764 42802
rect 10753 42756 10764 42773
rect 10810 42756 10878 42802
rect 10924 42756 10992 42802
rect 11038 42756 11106 42802
rect 11152 42756 11220 42802
rect 11266 42756 11334 42802
rect 11380 42756 11448 42802
rect 11494 42756 11562 42802
rect 11608 42756 11676 42802
rect 11722 42756 11790 42802
rect 11836 42756 12075 42802
rect 10753 42688 12075 42756
rect 10753 42642 10764 42688
rect 10810 42642 10878 42688
rect 10924 42642 10992 42688
rect 11038 42642 11106 42688
rect 11152 42642 11220 42688
rect 11266 42642 11334 42688
rect 11380 42642 11448 42688
rect 11494 42642 11562 42688
rect 11608 42642 11676 42688
rect 11722 42642 11790 42688
rect 11836 42642 12075 42688
rect 3608 42580 3684 42592
rect 3608 41280 3620 42580
rect 3672 41280 3684 42580
rect 10753 42574 12075 42642
rect 10753 42528 10764 42574
rect 10810 42528 10878 42574
rect 10924 42528 10992 42574
rect 11038 42528 11106 42574
rect 11152 42528 11220 42574
rect 11266 42528 11334 42574
rect 11380 42528 11448 42574
rect 11494 42528 11562 42574
rect 11608 42528 11676 42574
rect 11722 42528 11790 42574
rect 11836 42528 12075 42574
rect 10753 42460 12075 42528
rect 10753 42414 10764 42460
rect 10810 42414 10878 42460
rect 10924 42414 10992 42460
rect 11038 42414 11106 42460
rect 11152 42414 11220 42460
rect 11266 42414 11334 42460
rect 11380 42414 11448 42460
rect 11494 42414 11562 42460
rect 11608 42414 11676 42460
rect 11722 42414 11790 42460
rect 11836 42414 12075 42460
rect 10753 42346 12075 42414
rect 10753 42300 10764 42346
rect 10810 42300 10878 42346
rect 10924 42300 10992 42346
rect 11038 42300 11106 42346
rect 11152 42300 11220 42346
rect 11266 42300 11334 42346
rect 11380 42300 11448 42346
rect 11494 42300 11562 42346
rect 11608 42300 11676 42346
rect 11722 42300 11790 42346
rect 11836 42300 12075 42346
rect 10753 42289 12075 42300
rect 3608 41268 3684 41280
rect 11290 41612 11826 41625
rect 11290 41566 11303 41612
rect 11349 41566 11419 41612
rect 11465 41566 11535 41612
rect 11581 41566 11651 41612
rect 11697 41566 11767 41612
rect 11813 41566 11826 41612
rect 11290 41553 11826 41566
rect 11290 41496 11362 41553
rect 11290 41450 11303 41496
rect 11349 41450 11362 41496
rect 11754 41496 11826 41553
rect 11290 41380 11362 41450
rect 11290 41334 11303 41380
rect 11349 41334 11362 41380
rect 11290 41264 11362 41334
rect 11290 41218 11303 41264
rect 11349 41218 11362 41264
rect 11458 41444 11658 41457
rect 11458 41398 11471 41444
rect 11458 41316 11517 41398
rect 11458 41270 11471 41316
rect 11569 41398 11599 41444
rect 11645 41398 11658 41444
rect 11569 41316 11658 41398
rect 11569 41288 11599 41316
rect 11517 41270 11599 41288
rect 11645 41270 11658 41316
rect 11458 41257 11658 41270
rect 11754 41450 11767 41496
rect 11813 41450 11826 41496
rect 11754 41380 11826 41450
rect 11754 41334 11767 41380
rect 11813 41334 11826 41380
rect 11754 41264 11826 41334
rect 11290 41161 11362 41218
rect 11754 41218 11767 41264
rect 11813 41218 11826 41264
rect 11754 41161 11826 41218
rect 11290 41148 11826 41161
rect 11290 41102 11303 41148
rect 11349 41102 11419 41148
rect 11465 41102 11535 41148
rect 11581 41102 11651 41148
rect 11697 41102 11767 41148
rect 11813 41102 11826 41148
rect 11290 41089 11826 41102
rect 11290 41032 11362 41089
rect 11290 40986 11303 41032
rect 11349 40986 11362 41032
rect 11754 41032 11826 41089
rect 11290 40916 11362 40986
rect 11290 40870 11303 40916
rect 11349 40870 11362 40916
rect 11290 40805 11362 40870
rect 11137 40800 11362 40805
rect 11137 40793 11303 40800
rect 1836 40700 3680 40712
rect 1836 40648 1848 40700
rect 3668 40648 3680 40700
rect 1836 40636 3680 40648
rect 11137 40637 11149 40793
rect 11201 40754 11303 40793
rect 11349 40754 11362 40800
rect 11458 40980 11658 40993
rect 11458 40934 11471 40980
rect 11517 40971 11599 40980
rect 11517 40934 11532 40971
rect 11458 40852 11532 40934
rect 11458 40806 11471 40852
rect 11517 40815 11532 40852
rect 11584 40934 11599 40971
rect 11645 40934 11658 40980
rect 11584 40852 11658 40934
rect 11584 40815 11599 40852
rect 11517 40806 11599 40815
rect 11645 40806 11658 40852
rect 11458 40793 11658 40806
rect 11754 40986 11767 41032
rect 11813 40986 11826 41032
rect 11754 40916 11826 40986
rect 11754 40870 11767 40916
rect 11813 40870 11826 40916
rect 11754 40800 11826 40870
rect 11201 40697 11362 40754
rect 11754 40754 11767 40800
rect 11813 40754 11826 40800
rect 11754 40697 11826 40754
rect 12064 40717 12075 42289
rect 12121 43161 12182 43207
rect 14484 43161 14592 43207
rect 12121 42821 14592 43161
rect 12121 42775 12519 42821
rect 13045 42775 13659 42821
rect 14185 42775 14592 42821
rect 12121 42764 14592 42775
rect 12121 42128 12332 42764
rect 12392 42693 13172 42704
rect 12392 42647 12403 42693
rect 12449 42647 13115 42693
rect 13161 42647 13172 42693
rect 12392 42581 13172 42647
rect 12392 42535 12403 42581
rect 12449 42535 13115 42581
rect 13161 42535 13172 42581
rect 12392 42498 13172 42535
rect 12392 42469 13108 42498
rect 13160 42469 13172 42498
rect 12392 42423 12403 42469
rect 12449 42423 13108 42469
rect 13161 42423 13172 42469
rect 12392 42357 13108 42423
rect 13160 42357 13172 42423
rect 12392 42311 12403 42357
rect 12449 42342 13108 42357
rect 12449 42311 13115 42342
rect 13161 42311 13172 42357
rect 12392 42245 13172 42311
rect 12392 42199 12403 42245
rect 12449 42199 13115 42245
rect 13161 42199 13172 42245
rect 12392 42188 13172 42199
rect 13272 42128 13472 42764
rect 13532 42693 14312 42704
rect 13532 42647 13543 42693
rect 13589 42647 14255 42693
rect 14301 42647 14312 42693
rect 13532 42581 14312 42647
rect 13532 42535 13543 42581
rect 13589 42535 14255 42581
rect 14301 42535 14312 42581
rect 13532 42498 14312 42535
rect 13532 42469 13544 42498
rect 13596 42469 14312 42498
rect 13532 42423 13543 42469
rect 13596 42423 14255 42469
rect 14301 42423 14312 42469
rect 13532 42357 13544 42423
rect 13596 42357 14312 42423
rect 13532 42311 13543 42357
rect 13596 42342 14255 42357
rect 13589 42311 14255 42342
rect 14301 42311 14312 42357
rect 13532 42245 14312 42311
rect 13532 42199 13543 42245
rect 13589 42199 14255 42245
rect 14301 42199 14312 42245
rect 13532 42188 14312 42199
rect 12121 42117 13082 42128
rect 12121 42071 12519 42117
rect 13045 42071 13082 42117
rect 12121 41853 13082 42071
rect 12121 41807 12519 41853
rect 13045 41807 13082 41853
rect 12121 41796 13082 41807
rect 13272 42117 14222 42128
rect 13272 42071 13659 42117
rect 14185 42071 14222 42117
rect 13272 41853 14222 42071
rect 13272 41807 13659 41853
rect 14185 41807 14222 41853
rect 13272 41796 14222 41807
rect 12121 41160 12332 41796
rect 12392 41725 13172 41736
rect 12392 41679 12403 41725
rect 12449 41679 13115 41725
rect 13161 41679 13172 41725
rect 12392 41613 13172 41679
rect 12392 41567 12403 41613
rect 12449 41571 13115 41613
rect 12449 41567 13108 41571
rect 13161 41567 13172 41613
rect 12392 41501 13108 41567
rect 13160 41501 13172 41567
rect 12392 41455 12403 41501
rect 12449 41455 13108 41501
rect 13161 41455 13172 41501
rect 12392 41415 13108 41455
rect 13160 41415 13172 41455
rect 12392 41389 13172 41415
rect 12392 41343 12403 41389
rect 12449 41343 13115 41389
rect 13161 41343 13172 41389
rect 12392 41277 13172 41343
rect 12392 41231 12403 41277
rect 12449 41231 13115 41277
rect 13161 41231 13172 41277
rect 12392 41220 13172 41231
rect 13272 41160 13472 41796
rect 13532 41725 14312 41736
rect 13532 41679 13543 41725
rect 13589 41679 14255 41725
rect 14301 41679 14312 41725
rect 13532 41613 14312 41679
rect 13532 41567 13543 41613
rect 13589 41571 14255 41613
rect 13596 41567 14255 41571
rect 14301 41567 14312 41613
rect 13532 41501 13544 41567
rect 13596 41501 14312 41567
rect 13532 41455 13543 41501
rect 13596 41455 14255 41501
rect 14301 41455 14312 41501
rect 13532 41415 13544 41455
rect 13596 41415 14312 41455
rect 13532 41389 14312 41415
rect 13532 41343 13543 41389
rect 13589 41343 14255 41389
rect 14301 41343 14312 41389
rect 13532 41277 14312 41343
rect 13532 41231 13543 41277
rect 13589 41231 14255 41277
rect 14301 41231 14312 41277
rect 13532 41220 14312 41231
rect 14581 41224 14592 42764
rect 14547 41160 14592 41224
rect 12121 41149 14592 41160
rect 12121 41103 12519 41149
rect 13045 41103 13659 41149
rect 14185 41103 14592 41149
rect 12121 40763 14592 41103
rect 12121 40717 12182 40763
rect 14484 40717 14592 40763
rect 14638 42764 14745 43207
rect 14638 41224 14649 42764
rect 14638 41160 14703 41224
rect 14638 40717 14745 41160
rect 12064 40706 14745 40717
rect 11201 40684 11826 40697
rect 11201 40638 11303 40684
rect 11349 40638 11419 40684
rect 11465 40638 11535 40684
rect 11581 40638 11651 40684
rect 11697 40638 11767 40684
rect 11813 40638 11826 40684
rect 11201 40637 11826 40638
rect 11137 40625 11826 40637
rect 14058 40468 14134 40480
rect 14058 40376 14070 40468
rect 1913 40364 14070 40376
rect 1913 40312 1925 40364
rect 2081 40312 4849 40364
rect 5005 40312 7065 40364
rect 7221 40312 10796 40364
rect 10952 40312 14070 40364
rect 14122 40312 14134 40468
rect 1913 40300 14134 40312
rect 1596 40228 5746 40240
rect 1596 40176 1608 40228
rect 1764 40176 5578 40228
rect 5734 40176 5746 40228
rect 1596 40164 5746 40176
rect 11416 40228 13842 40240
rect 11416 40176 11428 40228
rect 11584 40176 13674 40228
rect 13830 40176 13842 40228
rect 11416 40164 13842 40176
rect 10644 40092 13988 40104
rect 10644 40040 10656 40092
rect 10812 40040 11996 40092
rect 12152 40040 13820 40092
rect 13976 40040 13988 40092
rect 10644 40028 13988 40040
rect 184 39936 954 39948
rect 184 39884 202 39936
rect 566 39884 954 39936
rect 184 39880 954 39884
rect 2433 39944 4485 39956
rect 2433 39892 2445 39944
rect 4473 39892 4485 39944
rect 2433 39880 4485 39892
rect 7888 39944 9732 39956
rect 7888 39892 7900 39944
rect 9720 39892 9732 39944
rect 7888 39880 9732 39892
rect 12772 39944 13784 39956
rect 12772 39892 12784 39944
rect 13772 39892 13784 39944
rect 12772 39880 13784 39892
rect 190 39872 578 39880
rect 14323 39709 14523 40706
rect 14193 39509 14523 39709
rect 1771 39418 1847 39430
rect 1771 38846 1783 39418
rect 1835 38846 1847 39418
rect 1771 38834 1847 38846
rect 5083 39418 5159 39430
rect 5083 38846 5095 39418
rect 5147 38846 5159 39418
rect 5083 38834 5159 38846
rect 6049 39418 6125 39430
rect 6049 38430 6061 39418
rect 6113 38430 6125 39418
rect 7015 39418 7091 39430
rect 6306 38687 6382 39089
rect 7015 38846 7027 39418
rect 7079 38846 7091 39418
rect 7015 38834 7091 38846
rect 10327 39418 10403 39430
rect 6306 38507 6504 38687
rect 6049 38418 6125 38430
rect 10327 38430 10339 39418
rect 10391 38430 10403 39418
rect 11200 39418 11276 39430
rect 10644 38676 10720 38688
rect 10644 38520 10656 38676
rect 10708 38520 10720 38676
rect 10644 38508 10720 38520
rect 10888 38676 10964 38688
rect 10888 38520 10900 38676
rect 10952 38520 10964 38676
rect 10888 38508 10964 38520
rect 10327 38418 10403 38430
rect 11200 38430 11212 39418
rect 11264 38430 11276 39418
rect 11200 38418 11276 38430
rect 8293 38318 8369 38330
rect 8293 38162 8305 38318
rect 8357 38162 8369 38318
rect 0 36480 58 37780
rect 110 36480 122 37780
rect 805 38142 881 38154
rect 805 37154 817 38142
rect 869 37154 881 38142
rect 3427 38142 3503 38154
rect 2707 37569 2783 37581
rect 2707 37413 2719 37569
rect 2771 37413 2783 37569
rect 2707 37401 2783 37413
rect 3195 37569 3271 37581
rect 3195 37413 3207 37569
rect 3259 37413 3271 37569
rect 3195 37401 3271 37413
rect 805 37142 881 37154
rect 3427 37154 3439 38142
rect 3491 37154 3503 38142
rect 6049 38142 6125 38154
rect 8293 38150 8369 38162
rect 11520 38315 11596 38327
rect 11520 38159 11532 38315
rect 11584 38159 11596 38315
rect 3659 37569 3735 37581
rect 3659 37413 3671 37569
rect 3723 37413 3735 37569
rect 3659 37401 3735 37413
rect 4147 37569 4223 37581
rect 4147 37413 4159 37569
rect 4211 37413 4223 37569
rect 4147 37401 4223 37413
rect 3427 37142 3503 37154
rect 6049 37154 6061 38142
rect 6113 37154 6125 38142
rect 8671 38142 8747 38154
rect 11520 38147 11596 38159
rect 13303 38307 13379 38319
rect 13303 38151 13315 38307
rect 13367 38151 13379 38307
rect 8439 37569 8515 37581
rect 8439 37413 8451 37569
rect 8503 37413 8515 37569
rect 8439 37401 8515 37413
rect 6049 37142 6125 37154
rect 8671 37154 8683 38142
rect 8735 37154 8747 38142
rect 13303 38139 13379 38151
rect 14193 38150 14393 39509
rect 13919 37910 14393 38150
rect 13439 37653 13515 37665
rect 8895 37569 8971 37581
rect 8895 37413 8907 37569
rect 8959 37413 8971 37569
rect 13439 37497 13451 37653
rect 13503 37497 13515 37653
rect 13439 37485 13515 37497
rect 8895 37401 8971 37413
rect 8671 37142 8747 37154
rect 10331 37198 11551 37210
rect 10331 37146 10343 37198
rect 11539 37146 11551 37198
rect 10331 37134 11551 37146
rect 0 9276 122 36480
rect 8439 36632 8515 36644
rect 8439 36476 8451 36632
rect 8503 36540 8515 36632
rect 8503 36528 13242 36540
rect 8503 36476 13074 36528
rect 13230 36476 13242 36528
rect 8439 36464 13242 36476
rect 8293 36392 13102 36404
rect 8293 36340 8305 36392
rect 8461 36340 12934 36392
rect 13090 36340 13102 36392
rect 8293 36328 13102 36340
rect 2066 36256 2469 36268
rect 2066 36204 2088 36256
rect 2452 36204 2469 36256
rect 2066 36192 2469 36204
rect 4461 36256 9150 36268
rect 4461 36204 4473 36256
rect 4629 36204 5822 36256
rect 5978 36204 8982 36256
rect 9138 36204 9150 36256
rect 4461 36192 9150 36204
rect 1822 36120 3271 36132
rect 1822 36068 1834 36120
rect 1990 36068 3103 36120
rect 3259 36068 3271 36120
rect 1822 36056 3271 36068
rect 3659 36120 9010 36132
rect 3659 36068 3671 36120
rect 3827 36068 6066 36120
rect 6222 36068 8842 36120
rect 8998 36068 9010 36120
rect 3659 36056 9010 36068
rect 2482 35984 12686 35996
rect 2482 35932 2494 35984
rect 2650 35932 5406 35984
rect 5562 35932 9502 35984
rect 9658 35932 12518 35984
rect 12674 35932 12686 35984
rect 2482 35920 12686 35932
rect 1310 35848 13754 35860
rect 1310 35796 1322 35848
rect 1478 35796 6578 35848
rect 6734 35796 8330 35848
rect 8486 35796 13586 35848
rect 13742 35796 13754 35848
rect 1310 35784 13754 35796
rect 3386 35712 13515 35724
rect 3386 35660 3398 35712
rect 3554 35660 4502 35712
rect 4658 35660 10406 35712
rect 10562 35660 11510 35712
rect 11666 35660 13347 35712
rect 13503 35660 13515 35712
rect 3386 35648 13515 35660
rect 486 35576 562 35588
rect 486 33756 498 35576
rect 550 33756 562 35576
rect 724 35576 800 35588
rect 724 34172 736 35576
rect 788 34172 800 35576
rect 724 34160 800 34172
rect 3092 35576 3168 35588
rect 3092 34172 3104 35576
rect 3156 34172 3168 35576
rect 3092 34160 3168 34172
rect 3990 35576 4066 35588
rect 1822 34065 1898 34077
rect 1822 33909 1834 34065
rect 1886 33909 1898 34065
rect 1822 33897 1898 33909
rect 2066 34065 2142 34077
rect 2066 33909 2078 34065
rect 2130 33909 2142 34065
rect 2066 33897 2142 33909
rect 2482 34065 2558 34077
rect 2482 33909 2494 34065
rect 2546 33909 2558 34065
rect 2482 33897 2558 33909
rect 486 33744 562 33756
rect 486 33481 562 33493
rect 486 29685 498 33481
rect 550 29685 562 33481
rect 3990 32924 4002 35576
rect 4054 32924 4066 35576
rect 4888 35576 4964 35588
rect 4888 34172 4900 35576
rect 4952 34172 4964 35576
rect 8567 35576 8747 35588
rect 8567 35524 8579 35576
rect 8735 35524 8747 35576
rect 8567 35512 8747 35524
rect 10100 35576 10176 35588
rect 4888 34160 4964 34172
rect 10100 34172 10112 35576
rect 10164 34172 10176 35576
rect 10100 34160 10176 34172
rect 10998 35576 11074 35588
rect 5498 34065 5574 34077
rect 5498 33909 5510 34065
rect 5562 33909 5574 34065
rect 5498 33897 5574 33909
rect 5914 34065 5990 34077
rect 5914 33909 5926 34065
rect 5978 33909 5990 34065
rect 5914 33897 5990 33909
rect 6158 34065 6234 34077
rect 6158 33909 6170 34065
rect 6222 33909 6234 34065
rect 6158 33897 6234 33909
rect 8830 34065 8906 34077
rect 8830 33909 8842 34065
rect 8894 33909 8906 34065
rect 8830 33897 8906 33909
rect 9074 34065 9150 34077
rect 9074 33909 9086 34065
rect 9138 33909 9150 34065
rect 9074 33897 9150 33909
rect 9490 34065 9566 34077
rect 9490 33909 9502 34065
rect 9554 33909 9566 34065
rect 9490 33897 9566 33909
rect 3990 32912 4066 32924
rect 10998 32924 11010 35576
rect 11062 32924 11074 35576
rect 11896 35576 11972 35588
rect 11896 34172 11908 35576
rect 11960 34172 11972 35576
rect 13919 35520 14119 37910
rect 14942 37780 15064 50880
rect 14942 36480 14954 37780
rect 15006 36480 15064 37780
rect 11896 34160 11972 34172
rect 12506 34065 12582 34077
rect 12506 33909 12518 34065
rect 12570 33909 12582 34065
rect 12506 33897 12582 33909
rect 12922 34065 12998 34077
rect 12922 33909 12934 34065
rect 12986 33909 12998 34065
rect 12922 33897 12998 33909
rect 13166 34065 13242 34077
rect 13166 33909 13178 34065
rect 13230 33909 13242 34065
rect 13166 33897 13242 33909
rect 10998 32912 11074 32924
rect 14502 33481 14578 33493
rect 3990 32455 4066 32467
rect 968 32320 1044 32332
rect 968 30084 980 32320
rect 1032 30084 1044 32320
rect 2360 32320 2436 32332
rect 968 30072 1044 30084
rect 1456 30308 1532 30320
rect 1456 29944 1468 30308
rect 1520 29944 1532 30308
rect 1456 29932 1532 29944
rect 1700 30308 1776 30320
rect 1700 29944 1712 30308
rect 1764 29944 1776 30308
rect 2360 30084 2372 32320
rect 2424 30084 2436 32320
rect 2360 30072 2436 30084
rect 2776 32320 2852 32332
rect 2776 30084 2788 32320
rect 2840 30084 2852 32320
rect 3264 32320 3340 32332
rect 3264 30708 3276 32320
rect 3328 30708 3340 32320
rect 3264 30696 3340 30708
rect 3752 32270 3828 32282
rect 3752 30658 3764 32270
rect 3816 30658 3828 32270
rect 3752 30646 3828 30658
rect 3990 30635 4002 32455
rect 4054 30635 4066 32455
rect 10998 32455 11074 32467
rect 4716 32320 4792 32332
rect 4228 32270 4304 32282
rect 4228 30658 4240 32270
rect 4292 30658 4304 32270
rect 4716 30708 4728 32320
rect 4780 30708 4792 32320
rect 4716 30696 4792 30708
rect 5204 32320 5280 32332
rect 5204 30708 5216 32320
rect 5268 30708 5280 32320
rect 5204 30696 5280 30708
rect 5620 32320 5696 32332
rect 5620 30708 5632 32320
rect 5684 30708 5696 32320
rect 5620 30696 5696 30708
rect 7012 32320 7088 32332
rect 4228 30646 4304 30658
rect 3990 30623 4066 30635
rect 3020 30488 3096 30500
rect 3020 30124 3032 30488
rect 3084 30124 3096 30488
rect 4472 30488 4548 30500
rect 3020 30112 3096 30124
rect 3508 30308 3584 30320
rect 2776 30072 2852 30084
rect 1700 29932 1776 29944
rect 3508 29944 3520 30308
rect 3572 29944 3584 30308
rect 4472 30124 4484 30488
rect 4536 30124 4548 30488
rect 4472 30112 4548 30124
rect 4960 30308 5036 30320
rect 3508 29932 3584 29944
rect 4960 29944 4972 30308
rect 5024 29944 5036 30308
rect 4960 29932 5036 29944
rect 6524 30308 6600 30320
rect 6524 29944 6536 30308
rect 6588 29944 6600 30308
rect 6524 29932 6600 29944
rect 6768 30308 6844 30320
rect 6768 29944 6780 30308
rect 6832 29944 6844 30308
rect 7012 30084 7024 32320
rect 7076 30084 7088 32320
rect 7012 30072 7088 30084
rect 7976 32320 8052 32332
rect 7976 30084 7988 32320
rect 8040 30084 8052 32320
rect 9368 32320 9444 32332
rect 9368 30708 9380 32320
rect 9432 30708 9444 32320
rect 9368 30696 9444 30708
rect 9784 32320 9860 32332
rect 9784 30708 9796 32320
rect 9848 30708 9860 32320
rect 9784 30696 9860 30708
rect 10272 32320 10348 32332
rect 10272 30708 10284 32320
rect 10336 30708 10348 32320
rect 10272 30696 10348 30708
rect 10760 32270 10836 32282
rect 10760 30658 10772 32270
rect 10824 30658 10836 32270
rect 10760 30646 10836 30658
rect 10998 30635 11010 32455
rect 11062 30635 11074 32455
rect 11724 32320 11800 32332
rect 11236 32270 11312 32282
rect 11236 30658 11248 32270
rect 11300 30658 11312 32270
rect 11724 30708 11736 32320
rect 11788 30708 11800 32320
rect 11724 30696 11800 30708
rect 12212 32320 12288 32332
rect 11236 30646 11312 30658
rect 10998 30623 11074 30635
rect 10516 30488 10592 30500
rect 7976 30072 8052 30084
rect 8464 30308 8540 30320
rect 6768 29932 6844 29944
rect 8464 29944 8476 30308
rect 8528 29944 8540 30308
rect 8464 29932 8540 29944
rect 8708 30308 8784 30320
rect 8708 29944 8720 30308
rect 8772 29944 8784 30308
rect 8708 29932 8784 29944
rect 10028 30308 10104 30320
rect 10028 29944 10040 30308
rect 10092 29944 10104 30308
rect 10516 30124 10528 30488
rect 10580 30124 10592 30488
rect 11968 30488 12044 30500
rect 10516 30112 10592 30124
rect 11480 30308 11556 30320
rect 10028 29932 10104 29944
rect 11480 29944 11492 30308
rect 11544 29944 11556 30308
rect 11968 30124 11980 30488
rect 12032 30124 12044 30488
rect 11968 30112 12044 30124
rect 12212 30084 12224 32320
rect 12276 30084 12288 32320
rect 12212 30072 12288 30084
rect 12628 32320 12704 32332
rect 12628 30084 12640 32320
rect 12692 30084 12704 32320
rect 14020 32320 14096 32332
rect 12628 30072 12704 30084
rect 13532 30308 13608 30320
rect 11480 29932 11556 29944
rect 13532 29944 13544 30308
rect 13596 29944 13608 30308
rect 13532 29932 13608 29944
rect 13776 30308 13852 30320
rect 13776 29944 13788 30308
rect 13840 29944 13852 30308
rect 14020 30084 14032 32320
rect 14084 30084 14096 32320
rect 14020 30072 14096 30084
rect 13776 29932 13852 29944
rect 486 29673 562 29685
rect 2000 29737 3324 29749
rect 2000 29685 2012 29737
rect 3312 29685 3324 29737
rect 2000 29673 3324 29685
rect 11937 29737 13261 29749
rect 11937 29685 11949 29737
rect 13249 29685 13261 29737
rect 11937 29673 13261 29685
rect 14502 29685 14514 33481
rect 14566 29685 14578 33481
rect 14502 29673 14578 29685
rect 1367 29447 6612 29471
rect 1367 29395 1379 29447
rect 1535 29395 6444 29447
rect 6600 29395 6612 29447
rect 1367 29371 6612 29395
rect 8696 29447 13699 29471
rect 8696 29395 8708 29447
rect 8864 29395 13531 29447
rect 13687 29395 13699 29447
rect 8696 29371 13699 29395
rect 1547 29267 6856 29291
rect 1547 29215 1559 29267
rect 1715 29215 6688 29267
rect 6844 29215 6856 29267
rect 1547 29191 6856 29215
rect 8452 29267 13519 29291
rect 8452 29215 8464 29267
rect 8620 29215 13351 29267
rect 13507 29215 13519 29267
rect 8452 29191 13519 29215
rect 2340 29060 3888 29111
rect 2340 29008 3508 29060
rect 3664 29008 3888 29060
rect 2340 28949 3888 29008
rect 2340 26120 2502 28949
rect 3726 26120 3888 28949
rect 4112 29099 4274 29111
rect 4112 28943 4167 29099
rect 4219 28943 4274 29099
rect 4112 26120 4274 28943
rect 4960 29099 5648 29111
rect 4960 28943 4972 29099
rect 5024 28949 5648 29099
rect 5024 28943 5036 28949
rect 4960 28931 5036 28943
rect 5486 26120 5648 28949
rect 5872 29099 7420 29111
rect 5872 28943 5926 29099
rect 5978 28949 7420 29099
rect 5978 28943 6034 28949
rect 5872 26120 6034 28943
rect 7258 26120 7420 28949
rect 7646 29099 9194 29111
rect 7646 28949 9088 29099
rect 7646 26120 7808 28949
rect 9032 28943 9088 28949
rect 9140 28943 9194 29099
rect 9032 26120 9194 28943
rect 9418 29099 10106 29111
rect 9418 28949 10042 29099
rect 9418 26120 9580 28949
rect 10030 28943 10042 28949
rect 10094 28943 10106 29099
rect 10030 28931 10106 28943
rect 10792 29099 10954 29111
rect 10792 28943 10847 29099
rect 10899 28943 10954 29099
rect 10792 26120 10954 28943
rect 11178 29060 12726 29111
rect 11178 29008 11402 29060
rect 11558 29008 12726 29060
rect 11178 28949 12726 29008
rect 11178 26120 11340 28949
rect 12564 26120 12726 28949
rect 14942 9276 15064 36480
rect 0 9265 832 9276
rect 0 9219 279 9265
rect 325 9219 403 9265
rect 449 9219 527 9265
rect 573 9219 651 9265
rect 697 9219 775 9265
rect 821 9219 832 9265
rect 0 9141 832 9219
rect 0 9095 279 9141
rect 325 9095 403 9141
rect 449 9095 527 9141
rect 573 9095 651 9141
rect 697 9095 775 9141
rect 821 9095 832 9141
rect 0 9017 832 9095
rect 0 8971 279 9017
rect 325 8971 403 9017
rect 449 8971 527 9017
rect 573 8971 651 9017
rect 697 8971 775 9017
rect 821 8971 832 9017
rect 0 8893 832 8971
rect 0 8847 279 8893
rect 325 8847 403 8893
rect 449 8847 527 8893
rect 573 8847 651 8893
rect 697 8847 775 8893
rect 821 8847 832 8893
rect 0 8769 832 8847
rect 0 8723 279 8769
rect 325 8723 403 8769
rect 449 8723 527 8769
rect 573 8723 651 8769
rect 697 8723 775 8769
rect 821 8723 832 8769
rect 0 8645 832 8723
rect 0 8599 279 8645
rect 325 8599 403 8645
rect 449 8599 527 8645
rect 573 8599 651 8645
rect 697 8599 775 8645
rect 821 8599 832 8645
rect 0 8521 832 8599
rect 0 8475 279 8521
rect 325 8475 403 8521
rect 449 8475 527 8521
rect 573 8475 651 8521
rect 697 8475 775 8521
rect 821 8475 832 8521
rect 0 8397 832 8475
rect 0 8351 279 8397
rect 325 8351 403 8397
rect 449 8351 527 8397
rect 573 8351 651 8397
rect 697 8351 775 8397
rect 821 8351 832 8397
rect 0 8273 832 8351
rect 0 8227 279 8273
rect 325 8227 403 8273
rect 449 8227 527 8273
rect 573 8227 651 8273
rect 697 8227 775 8273
rect 821 8227 832 8273
rect 0 8149 832 8227
rect 0 8103 279 8149
rect 325 8103 403 8149
rect 449 8103 527 8149
rect 573 8103 651 8149
rect 697 8103 775 8149
rect 821 8103 832 8149
rect 0 8025 832 8103
rect 0 7979 279 8025
rect 325 7979 403 8025
rect 449 7979 527 8025
rect 573 7979 651 8025
rect 697 7979 775 8025
rect 821 7979 832 8025
rect 0 7901 832 7979
rect 0 7855 279 7901
rect 325 7855 403 7901
rect 449 7855 527 7901
rect 573 7855 651 7901
rect 697 7855 775 7901
rect 821 7855 832 7901
rect 0 7777 832 7855
rect 0 7731 279 7777
rect 325 7731 403 7777
rect 449 7731 527 7777
rect 573 7731 651 7777
rect 697 7731 775 7777
rect 821 7731 832 7777
rect 0 7653 832 7731
rect 0 7607 279 7653
rect 325 7607 403 7653
rect 449 7607 527 7653
rect 573 7607 651 7653
rect 697 7607 775 7653
rect 821 7607 832 7653
rect 0 7529 832 7607
rect 0 7483 279 7529
rect 325 7483 403 7529
rect 449 7483 527 7529
rect 573 7483 651 7529
rect 697 7483 775 7529
rect 821 7483 832 7529
rect 0 7405 832 7483
rect 0 7359 279 7405
rect 325 7359 403 7405
rect 449 7359 527 7405
rect 573 7359 651 7405
rect 697 7359 775 7405
rect 821 7359 832 7405
rect 0 7281 832 7359
rect 0 7235 279 7281
rect 325 7235 403 7281
rect 449 7235 527 7281
rect 573 7235 651 7281
rect 697 7235 775 7281
rect 821 7235 832 7281
rect 0 7157 832 7235
rect 0 7111 279 7157
rect 325 7111 403 7157
rect 449 7111 527 7157
rect 573 7111 651 7157
rect 697 7111 775 7157
rect 821 7111 832 7157
rect 0 7033 832 7111
rect 0 6987 279 7033
rect 325 6987 403 7033
rect 449 6987 527 7033
rect 573 6987 651 7033
rect 697 6987 775 7033
rect 821 6987 832 7033
rect 0 6909 832 6987
rect 0 6863 279 6909
rect 325 6863 403 6909
rect 449 6863 527 6909
rect 573 6863 651 6909
rect 697 6863 775 6909
rect 821 6863 832 6909
rect 0 6785 832 6863
rect 0 6739 279 6785
rect 325 6739 403 6785
rect 449 6739 527 6785
rect 573 6739 651 6785
rect 697 6739 775 6785
rect 821 6739 832 6785
rect 0 6661 832 6739
rect 0 6615 279 6661
rect 325 6615 403 6661
rect 449 6615 527 6661
rect 573 6615 651 6661
rect 697 6615 775 6661
rect 821 6615 832 6661
rect 0 6537 832 6615
rect 0 6491 279 6537
rect 325 6491 403 6537
rect 449 6491 527 6537
rect 573 6491 651 6537
rect 697 6491 775 6537
rect 821 6491 832 6537
rect 0 6413 832 6491
rect 0 6367 279 6413
rect 325 6367 403 6413
rect 449 6367 527 6413
rect 573 6367 651 6413
rect 697 6367 775 6413
rect 821 6367 832 6413
rect 0 6289 832 6367
rect 0 6243 279 6289
rect 325 6243 403 6289
rect 449 6243 527 6289
rect 573 6243 651 6289
rect 697 6243 775 6289
rect 821 6243 832 6289
rect 0 6165 832 6243
rect 0 6119 279 6165
rect 325 6119 403 6165
rect 449 6119 527 6165
rect 573 6119 651 6165
rect 697 6119 775 6165
rect 821 6119 832 6165
rect 0 6041 832 6119
rect 0 5995 279 6041
rect 325 5995 403 6041
rect 449 5995 527 6041
rect 573 5995 651 6041
rect 697 5995 775 6041
rect 821 5995 832 6041
rect 0 5917 832 5995
rect 0 5871 279 5917
rect 325 5871 403 5917
rect 449 5871 527 5917
rect 573 5871 651 5917
rect 697 5871 775 5917
rect 821 5871 832 5917
rect 0 5793 832 5871
rect 0 5747 279 5793
rect 325 5747 403 5793
rect 449 5747 527 5793
rect 573 5747 651 5793
rect 697 5747 775 5793
rect 821 5747 832 5793
rect 0 5669 832 5747
rect 0 5623 279 5669
rect 325 5623 403 5669
rect 449 5623 527 5669
rect 573 5623 651 5669
rect 697 5623 775 5669
rect 821 5623 832 5669
rect 0 5545 832 5623
rect 0 5499 279 5545
rect 325 5499 403 5545
rect 449 5499 527 5545
rect 573 5499 651 5545
rect 697 5499 775 5545
rect 821 5499 832 5545
rect 0 5421 832 5499
rect 0 5375 279 5421
rect 325 5375 403 5421
rect 449 5375 527 5421
rect 573 5375 651 5421
rect 697 5375 775 5421
rect 821 5375 832 5421
rect 0 5297 832 5375
rect 0 5251 279 5297
rect 325 5251 403 5297
rect 449 5251 527 5297
rect 573 5251 651 5297
rect 697 5251 775 5297
rect 821 5251 832 5297
rect 0 5173 832 5251
rect 0 5127 279 5173
rect 325 5127 403 5173
rect 449 5127 527 5173
rect 573 5127 651 5173
rect 697 5127 775 5173
rect 821 5127 832 5173
rect 0 5049 832 5127
rect 0 5003 279 5049
rect 325 5003 403 5049
rect 449 5003 527 5049
rect 573 5003 651 5049
rect 697 5003 775 5049
rect 821 5003 832 5049
rect 0 4925 832 5003
rect 0 4879 279 4925
rect 325 4879 403 4925
rect 449 4879 527 4925
rect 573 4879 651 4925
rect 697 4879 775 4925
rect 821 4879 832 4925
rect 0 4801 832 4879
rect 0 4755 279 4801
rect 325 4755 403 4801
rect 449 4755 527 4801
rect 573 4755 651 4801
rect 697 4755 775 4801
rect 821 4755 832 4801
rect 0 4677 832 4755
rect 0 4631 279 4677
rect 325 4631 403 4677
rect 449 4631 527 4677
rect 573 4631 651 4677
rect 697 4631 775 4677
rect 821 4631 832 4677
rect 0 4553 832 4631
rect 0 4507 279 4553
rect 325 4507 403 4553
rect 449 4507 527 4553
rect 573 4507 651 4553
rect 697 4507 775 4553
rect 821 4507 832 4553
rect 0 4429 832 4507
rect 0 4383 279 4429
rect 325 4383 403 4429
rect 449 4383 527 4429
rect 573 4383 651 4429
rect 697 4383 775 4429
rect 821 4383 832 4429
rect 0 4305 832 4383
rect 0 4259 279 4305
rect 325 4259 403 4305
rect 449 4259 527 4305
rect 573 4259 651 4305
rect 697 4259 775 4305
rect 821 4259 832 4305
rect 0 4181 832 4259
rect 0 4135 279 4181
rect 325 4135 403 4181
rect 449 4135 527 4181
rect 573 4135 651 4181
rect 697 4135 775 4181
rect 821 4135 832 4181
rect 0 4057 832 4135
rect 0 4011 279 4057
rect 325 4011 403 4057
rect 449 4011 527 4057
rect 573 4011 651 4057
rect 697 4011 775 4057
rect 821 4011 832 4057
rect 0 3933 832 4011
rect 0 3887 279 3933
rect 325 3887 403 3933
rect 449 3887 527 3933
rect 573 3887 651 3933
rect 697 3887 775 3933
rect 821 3887 832 3933
rect 0 3809 832 3887
rect 0 3763 279 3809
rect 325 3763 403 3809
rect 449 3763 527 3809
rect 573 3763 651 3809
rect 697 3763 775 3809
rect 821 3763 832 3809
rect 0 3685 832 3763
rect 0 3639 279 3685
rect 325 3639 403 3685
rect 449 3639 527 3685
rect 573 3639 651 3685
rect 697 3639 775 3685
rect 821 3639 832 3685
rect 0 3561 832 3639
rect 0 3515 279 3561
rect 325 3515 403 3561
rect 449 3515 527 3561
rect 573 3515 651 3561
rect 697 3515 775 3561
rect 821 3515 832 3561
rect 0 3437 832 3515
rect 0 3391 279 3437
rect 325 3391 403 3437
rect 449 3391 527 3437
rect 573 3391 651 3437
rect 697 3391 775 3437
rect 821 3391 832 3437
rect 0 3313 832 3391
rect 0 3267 279 3313
rect 325 3267 403 3313
rect 449 3267 527 3313
rect 573 3267 651 3313
rect 697 3267 775 3313
rect 821 3267 832 3313
rect 0 3189 832 3267
rect 0 3143 279 3189
rect 325 3143 403 3189
rect 449 3143 527 3189
rect 573 3143 651 3189
rect 697 3143 775 3189
rect 821 3143 832 3189
rect 0 3065 832 3143
rect 0 3019 279 3065
rect 325 3019 403 3065
rect 449 3019 527 3065
rect 573 3019 651 3065
rect 697 3019 775 3065
rect 821 3019 832 3065
rect 0 2941 832 3019
rect 0 2895 279 2941
rect 325 2895 403 2941
rect 449 2895 527 2941
rect 573 2895 651 2941
rect 697 2895 775 2941
rect 821 2895 832 2941
rect 0 2817 832 2895
rect 0 2771 279 2817
rect 325 2771 403 2817
rect 449 2771 527 2817
rect 573 2771 651 2817
rect 697 2771 775 2817
rect 821 2771 832 2817
rect 0 2693 832 2771
rect 0 2647 279 2693
rect 325 2647 403 2693
rect 449 2647 527 2693
rect 573 2647 651 2693
rect 697 2647 775 2693
rect 821 2647 832 2693
rect 0 2569 832 2647
rect 0 2523 279 2569
rect 325 2523 403 2569
rect 449 2523 527 2569
rect 573 2523 651 2569
rect 697 2523 775 2569
rect 821 2523 832 2569
rect 0 2445 832 2523
rect 0 2399 279 2445
rect 325 2399 403 2445
rect 449 2399 527 2445
rect 573 2399 651 2445
rect 697 2399 775 2445
rect 821 2399 832 2445
rect 0 2321 832 2399
rect 0 2275 279 2321
rect 325 2275 403 2321
rect 449 2275 527 2321
rect 573 2275 651 2321
rect 697 2275 775 2321
rect 821 2275 832 2321
rect 0 2197 832 2275
rect 0 2151 279 2197
rect 325 2151 403 2197
rect 449 2151 527 2197
rect 573 2151 651 2197
rect 697 2151 775 2197
rect 821 2151 832 2197
rect 0 2073 832 2151
rect 0 2027 279 2073
rect 325 2027 403 2073
rect 449 2027 527 2073
rect 573 2027 651 2073
rect 697 2027 775 2073
rect 821 2027 832 2073
rect 0 1949 832 2027
rect 0 1903 279 1949
rect 325 1903 403 1949
rect 449 1903 527 1949
rect 573 1903 651 1949
rect 697 1903 775 1949
rect 821 1903 832 1949
rect 0 1825 832 1903
rect 0 1779 279 1825
rect 325 1779 403 1825
rect 449 1779 527 1825
rect 573 1779 651 1825
rect 697 1779 775 1825
rect 821 1779 832 1825
rect 0 1701 832 1779
rect 0 1655 279 1701
rect 325 1655 403 1701
rect 449 1655 527 1701
rect 573 1655 651 1701
rect 697 1655 775 1701
rect 821 1655 832 1701
rect 0 1577 832 1655
rect 0 1531 279 1577
rect 325 1531 403 1577
rect 449 1531 527 1577
rect 573 1531 651 1577
rect 697 1531 775 1577
rect 821 1531 832 1577
rect 0 1453 832 1531
rect 0 1407 279 1453
rect 325 1407 403 1453
rect 449 1407 527 1453
rect 573 1407 651 1453
rect 697 1407 775 1453
rect 821 1407 832 1453
rect 0 1329 832 1407
rect 0 1283 279 1329
rect 325 1283 403 1329
rect 449 1283 527 1329
rect 573 1283 651 1329
rect 697 1283 775 1329
rect 821 1283 832 1329
rect 0 1205 832 1283
rect 0 1159 279 1205
rect 325 1159 403 1205
rect 449 1159 527 1205
rect 573 1159 651 1205
rect 697 1159 775 1205
rect 821 1159 832 1205
rect 0 1081 832 1159
rect 0 1035 279 1081
rect 325 1035 403 1081
rect 449 1035 527 1081
rect 573 1035 651 1081
rect 697 1035 775 1081
rect 821 1035 832 1081
rect 0 957 832 1035
rect 0 911 279 957
rect 325 911 403 957
rect 449 911 527 957
rect 573 911 651 957
rect 697 911 775 957
rect 821 911 832 957
rect 0 833 832 911
rect 0 787 279 833
rect 325 787 403 833
rect 449 787 527 833
rect 573 787 651 833
rect 697 787 775 833
rect 821 787 832 833
rect 0 709 832 787
rect 0 663 279 709
rect 325 663 403 709
rect 449 663 527 709
rect 573 663 651 709
rect 697 663 775 709
rect 821 663 832 709
rect 0 496 832 663
rect 14214 9265 15064 9276
rect 14214 9219 14225 9265
rect 14271 9219 14349 9265
rect 14395 9219 14473 9265
rect 14519 9219 14597 9265
rect 14643 9219 14721 9265
rect 14767 9219 15064 9265
rect 14214 9141 15064 9219
rect 14214 9095 14225 9141
rect 14271 9095 14349 9141
rect 14395 9095 14473 9141
rect 14519 9095 14597 9141
rect 14643 9095 14721 9141
rect 14767 9095 15064 9141
rect 14214 9017 15064 9095
rect 14214 8971 14225 9017
rect 14271 8971 14349 9017
rect 14395 8971 14473 9017
rect 14519 8971 14597 9017
rect 14643 8971 14721 9017
rect 14767 8971 15064 9017
rect 14214 8893 15064 8971
rect 14214 8847 14225 8893
rect 14271 8847 14349 8893
rect 14395 8847 14473 8893
rect 14519 8847 14597 8893
rect 14643 8847 14721 8893
rect 14767 8847 15064 8893
rect 14214 8769 15064 8847
rect 14214 8723 14225 8769
rect 14271 8723 14349 8769
rect 14395 8723 14473 8769
rect 14519 8723 14597 8769
rect 14643 8723 14721 8769
rect 14767 8723 15064 8769
rect 14214 8645 15064 8723
rect 14214 8599 14225 8645
rect 14271 8599 14349 8645
rect 14395 8599 14473 8645
rect 14519 8599 14597 8645
rect 14643 8599 14721 8645
rect 14767 8599 15064 8645
rect 14214 8521 15064 8599
rect 14214 8475 14225 8521
rect 14271 8475 14349 8521
rect 14395 8475 14473 8521
rect 14519 8475 14597 8521
rect 14643 8475 14721 8521
rect 14767 8475 15064 8521
rect 14214 8397 15064 8475
rect 14214 8351 14225 8397
rect 14271 8351 14349 8397
rect 14395 8351 14473 8397
rect 14519 8351 14597 8397
rect 14643 8351 14721 8397
rect 14767 8351 15064 8397
rect 14214 8273 15064 8351
rect 14214 8227 14225 8273
rect 14271 8227 14349 8273
rect 14395 8227 14473 8273
rect 14519 8227 14597 8273
rect 14643 8227 14721 8273
rect 14767 8227 15064 8273
rect 14214 8149 15064 8227
rect 14214 8103 14225 8149
rect 14271 8103 14349 8149
rect 14395 8103 14473 8149
rect 14519 8103 14597 8149
rect 14643 8103 14721 8149
rect 14767 8103 15064 8149
rect 14214 8025 15064 8103
rect 14214 7979 14225 8025
rect 14271 7979 14349 8025
rect 14395 7979 14473 8025
rect 14519 7979 14597 8025
rect 14643 7979 14721 8025
rect 14767 7979 15064 8025
rect 14214 7901 15064 7979
rect 14214 7855 14225 7901
rect 14271 7855 14349 7901
rect 14395 7855 14473 7901
rect 14519 7855 14597 7901
rect 14643 7855 14721 7901
rect 14767 7855 15064 7901
rect 14214 7777 15064 7855
rect 14214 7731 14225 7777
rect 14271 7731 14349 7777
rect 14395 7731 14473 7777
rect 14519 7731 14597 7777
rect 14643 7731 14721 7777
rect 14767 7731 15064 7777
rect 14214 7653 15064 7731
rect 14214 7607 14225 7653
rect 14271 7607 14349 7653
rect 14395 7607 14473 7653
rect 14519 7607 14597 7653
rect 14643 7607 14721 7653
rect 14767 7607 15064 7653
rect 14214 7529 15064 7607
rect 14214 7483 14225 7529
rect 14271 7483 14349 7529
rect 14395 7483 14473 7529
rect 14519 7483 14597 7529
rect 14643 7483 14721 7529
rect 14767 7483 15064 7529
rect 14214 7405 15064 7483
rect 14214 7359 14225 7405
rect 14271 7359 14349 7405
rect 14395 7359 14473 7405
rect 14519 7359 14597 7405
rect 14643 7359 14721 7405
rect 14767 7359 15064 7405
rect 14214 7281 15064 7359
rect 14214 7235 14225 7281
rect 14271 7235 14349 7281
rect 14395 7235 14473 7281
rect 14519 7235 14597 7281
rect 14643 7235 14721 7281
rect 14767 7235 15064 7281
rect 14214 7157 15064 7235
rect 14214 7111 14225 7157
rect 14271 7111 14349 7157
rect 14395 7111 14473 7157
rect 14519 7111 14597 7157
rect 14643 7111 14721 7157
rect 14767 7111 15064 7157
rect 14214 7033 15064 7111
rect 14214 6987 14225 7033
rect 14271 6987 14349 7033
rect 14395 6987 14473 7033
rect 14519 6987 14597 7033
rect 14643 6987 14721 7033
rect 14767 6987 15064 7033
rect 14214 6909 15064 6987
rect 14214 6863 14225 6909
rect 14271 6863 14349 6909
rect 14395 6863 14473 6909
rect 14519 6863 14597 6909
rect 14643 6863 14721 6909
rect 14767 6863 15064 6909
rect 14214 6785 15064 6863
rect 14214 6739 14225 6785
rect 14271 6739 14349 6785
rect 14395 6739 14473 6785
rect 14519 6739 14597 6785
rect 14643 6739 14721 6785
rect 14767 6739 15064 6785
rect 14214 6661 15064 6739
rect 14214 6615 14225 6661
rect 14271 6615 14349 6661
rect 14395 6615 14473 6661
rect 14519 6615 14597 6661
rect 14643 6615 14721 6661
rect 14767 6615 15064 6661
rect 14214 6537 15064 6615
rect 14214 6491 14225 6537
rect 14271 6491 14349 6537
rect 14395 6491 14473 6537
rect 14519 6491 14597 6537
rect 14643 6491 14721 6537
rect 14767 6491 15064 6537
rect 14214 6413 15064 6491
rect 14214 6367 14225 6413
rect 14271 6367 14349 6413
rect 14395 6367 14473 6413
rect 14519 6367 14597 6413
rect 14643 6367 14721 6413
rect 14767 6367 15064 6413
rect 14214 6289 15064 6367
rect 14214 6243 14225 6289
rect 14271 6243 14349 6289
rect 14395 6243 14473 6289
rect 14519 6243 14597 6289
rect 14643 6243 14721 6289
rect 14767 6243 15064 6289
rect 14214 6165 15064 6243
rect 14214 6119 14225 6165
rect 14271 6119 14349 6165
rect 14395 6119 14473 6165
rect 14519 6119 14597 6165
rect 14643 6119 14721 6165
rect 14767 6119 15064 6165
rect 14214 6041 15064 6119
rect 14214 5995 14225 6041
rect 14271 5995 14349 6041
rect 14395 5995 14473 6041
rect 14519 5995 14597 6041
rect 14643 5995 14721 6041
rect 14767 5995 15064 6041
rect 14214 5917 15064 5995
rect 14214 5871 14225 5917
rect 14271 5871 14349 5917
rect 14395 5871 14473 5917
rect 14519 5871 14597 5917
rect 14643 5871 14721 5917
rect 14767 5871 15064 5917
rect 14214 5793 15064 5871
rect 14214 5747 14225 5793
rect 14271 5747 14349 5793
rect 14395 5747 14473 5793
rect 14519 5747 14597 5793
rect 14643 5747 14721 5793
rect 14767 5747 15064 5793
rect 14214 5669 15064 5747
rect 14214 5623 14225 5669
rect 14271 5623 14349 5669
rect 14395 5623 14473 5669
rect 14519 5623 14597 5669
rect 14643 5623 14721 5669
rect 14767 5623 15064 5669
rect 14214 5545 15064 5623
rect 14214 5499 14225 5545
rect 14271 5499 14349 5545
rect 14395 5499 14473 5545
rect 14519 5499 14597 5545
rect 14643 5499 14721 5545
rect 14767 5499 15064 5545
rect 14214 5421 15064 5499
rect 14214 5375 14225 5421
rect 14271 5375 14349 5421
rect 14395 5375 14473 5421
rect 14519 5375 14597 5421
rect 14643 5375 14721 5421
rect 14767 5375 15064 5421
rect 14214 5297 15064 5375
rect 14214 5251 14225 5297
rect 14271 5251 14349 5297
rect 14395 5251 14473 5297
rect 14519 5251 14597 5297
rect 14643 5251 14721 5297
rect 14767 5251 15064 5297
rect 14214 5173 15064 5251
rect 14214 5127 14225 5173
rect 14271 5127 14349 5173
rect 14395 5127 14473 5173
rect 14519 5127 14597 5173
rect 14643 5127 14721 5173
rect 14767 5127 15064 5173
rect 14214 5049 15064 5127
rect 14214 5003 14225 5049
rect 14271 5003 14349 5049
rect 14395 5003 14473 5049
rect 14519 5003 14597 5049
rect 14643 5003 14721 5049
rect 14767 5003 15064 5049
rect 14214 4925 15064 5003
rect 14214 4879 14225 4925
rect 14271 4879 14349 4925
rect 14395 4879 14473 4925
rect 14519 4879 14597 4925
rect 14643 4879 14721 4925
rect 14767 4879 15064 4925
rect 14214 4801 15064 4879
rect 14214 4755 14225 4801
rect 14271 4755 14349 4801
rect 14395 4755 14473 4801
rect 14519 4755 14597 4801
rect 14643 4755 14721 4801
rect 14767 4755 15064 4801
rect 14214 4677 15064 4755
rect 14214 4631 14225 4677
rect 14271 4631 14349 4677
rect 14395 4631 14473 4677
rect 14519 4631 14597 4677
rect 14643 4631 14721 4677
rect 14767 4631 15064 4677
rect 14214 4553 15064 4631
rect 14214 4507 14225 4553
rect 14271 4507 14349 4553
rect 14395 4507 14473 4553
rect 14519 4507 14597 4553
rect 14643 4507 14721 4553
rect 14767 4507 15064 4553
rect 14214 4429 15064 4507
rect 14214 4383 14225 4429
rect 14271 4383 14349 4429
rect 14395 4383 14473 4429
rect 14519 4383 14597 4429
rect 14643 4383 14721 4429
rect 14767 4383 15064 4429
rect 14214 4305 15064 4383
rect 14214 4259 14225 4305
rect 14271 4259 14349 4305
rect 14395 4259 14473 4305
rect 14519 4259 14597 4305
rect 14643 4259 14721 4305
rect 14767 4259 15064 4305
rect 14214 4181 15064 4259
rect 14214 4135 14225 4181
rect 14271 4135 14349 4181
rect 14395 4135 14473 4181
rect 14519 4135 14597 4181
rect 14643 4135 14721 4181
rect 14767 4135 15064 4181
rect 14214 4057 15064 4135
rect 14214 4011 14225 4057
rect 14271 4011 14349 4057
rect 14395 4011 14473 4057
rect 14519 4011 14597 4057
rect 14643 4011 14721 4057
rect 14767 4011 15064 4057
rect 14214 3933 15064 4011
rect 14214 3887 14225 3933
rect 14271 3887 14349 3933
rect 14395 3887 14473 3933
rect 14519 3887 14597 3933
rect 14643 3887 14721 3933
rect 14767 3887 15064 3933
rect 14214 3809 15064 3887
rect 14214 3763 14225 3809
rect 14271 3763 14349 3809
rect 14395 3763 14473 3809
rect 14519 3763 14597 3809
rect 14643 3763 14721 3809
rect 14767 3763 15064 3809
rect 14214 3685 15064 3763
rect 14214 3639 14225 3685
rect 14271 3639 14349 3685
rect 14395 3639 14473 3685
rect 14519 3639 14597 3685
rect 14643 3639 14721 3685
rect 14767 3639 15064 3685
rect 14214 3561 15064 3639
rect 14214 3515 14225 3561
rect 14271 3515 14349 3561
rect 14395 3515 14473 3561
rect 14519 3515 14597 3561
rect 14643 3515 14721 3561
rect 14767 3515 15064 3561
rect 14214 3437 15064 3515
rect 14214 3391 14225 3437
rect 14271 3391 14349 3437
rect 14395 3391 14473 3437
rect 14519 3391 14597 3437
rect 14643 3391 14721 3437
rect 14767 3391 15064 3437
rect 14214 3313 15064 3391
rect 14214 3267 14225 3313
rect 14271 3267 14349 3313
rect 14395 3267 14473 3313
rect 14519 3267 14597 3313
rect 14643 3267 14721 3313
rect 14767 3267 15064 3313
rect 14214 3189 15064 3267
rect 14214 3143 14225 3189
rect 14271 3143 14349 3189
rect 14395 3143 14473 3189
rect 14519 3143 14597 3189
rect 14643 3143 14721 3189
rect 14767 3143 15064 3189
rect 14214 3065 15064 3143
rect 14214 3019 14225 3065
rect 14271 3019 14349 3065
rect 14395 3019 14473 3065
rect 14519 3019 14597 3065
rect 14643 3019 14721 3065
rect 14767 3019 15064 3065
rect 14214 2941 15064 3019
rect 14214 2895 14225 2941
rect 14271 2895 14349 2941
rect 14395 2895 14473 2941
rect 14519 2895 14597 2941
rect 14643 2895 14721 2941
rect 14767 2895 15064 2941
rect 14214 2817 15064 2895
rect 14214 2771 14225 2817
rect 14271 2771 14349 2817
rect 14395 2771 14473 2817
rect 14519 2771 14597 2817
rect 14643 2771 14721 2817
rect 14767 2771 15064 2817
rect 14214 2693 15064 2771
rect 14214 2647 14225 2693
rect 14271 2647 14349 2693
rect 14395 2647 14473 2693
rect 14519 2647 14597 2693
rect 14643 2647 14721 2693
rect 14767 2647 15064 2693
rect 14214 2569 15064 2647
rect 14214 2523 14225 2569
rect 14271 2523 14349 2569
rect 14395 2523 14473 2569
rect 14519 2523 14597 2569
rect 14643 2523 14721 2569
rect 14767 2523 15064 2569
rect 14214 2445 15064 2523
rect 14214 2399 14225 2445
rect 14271 2399 14349 2445
rect 14395 2399 14473 2445
rect 14519 2399 14597 2445
rect 14643 2399 14721 2445
rect 14767 2399 15064 2445
rect 14214 2321 15064 2399
rect 14214 2275 14225 2321
rect 14271 2275 14349 2321
rect 14395 2275 14473 2321
rect 14519 2275 14597 2321
rect 14643 2275 14721 2321
rect 14767 2275 15064 2321
rect 14214 2197 15064 2275
rect 14214 2151 14225 2197
rect 14271 2151 14349 2197
rect 14395 2151 14473 2197
rect 14519 2151 14597 2197
rect 14643 2151 14721 2197
rect 14767 2151 15064 2197
rect 14214 2073 15064 2151
rect 14214 2027 14225 2073
rect 14271 2027 14349 2073
rect 14395 2027 14473 2073
rect 14519 2027 14597 2073
rect 14643 2027 14721 2073
rect 14767 2027 15064 2073
rect 14214 1949 15064 2027
rect 14214 1903 14225 1949
rect 14271 1903 14349 1949
rect 14395 1903 14473 1949
rect 14519 1903 14597 1949
rect 14643 1903 14721 1949
rect 14767 1903 15064 1949
rect 14214 1825 15064 1903
rect 14214 1779 14225 1825
rect 14271 1779 14349 1825
rect 14395 1779 14473 1825
rect 14519 1779 14597 1825
rect 14643 1779 14721 1825
rect 14767 1779 15064 1825
rect 14214 1701 15064 1779
rect 14214 1655 14225 1701
rect 14271 1655 14349 1701
rect 14395 1655 14473 1701
rect 14519 1655 14597 1701
rect 14643 1655 14721 1701
rect 14767 1655 15064 1701
rect 14214 1577 15064 1655
rect 14214 1531 14225 1577
rect 14271 1531 14349 1577
rect 14395 1531 14473 1577
rect 14519 1531 14597 1577
rect 14643 1531 14721 1577
rect 14767 1531 15064 1577
rect 14214 1453 15064 1531
rect 14214 1407 14225 1453
rect 14271 1407 14349 1453
rect 14395 1407 14473 1453
rect 14519 1407 14597 1453
rect 14643 1407 14721 1453
rect 14767 1407 15064 1453
rect 14214 1329 15064 1407
rect 14214 1283 14225 1329
rect 14271 1283 14349 1329
rect 14395 1283 14473 1329
rect 14519 1283 14597 1329
rect 14643 1283 14721 1329
rect 14767 1283 15064 1329
rect 14214 1205 15064 1283
rect 14214 1159 14225 1205
rect 14271 1159 14349 1205
rect 14395 1159 14473 1205
rect 14519 1159 14597 1205
rect 14643 1159 14721 1205
rect 14767 1159 15064 1205
rect 14214 1081 15064 1159
rect 14214 1035 14225 1081
rect 14271 1035 14349 1081
rect 14395 1035 14473 1081
rect 14519 1035 14597 1081
rect 14643 1035 14721 1081
rect 14767 1035 15064 1081
rect 14214 957 15064 1035
rect 14214 911 14225 957
rect 14271 911 14349 957
rect 14395 911 14473 957
rect 14519 911 14597 957
rect 14643 911 14721 957
rect 14767 911 15064 957
rect 14214 833 15064 911
rect 14214 787 14225 833
rect 14271 787 14349 833
rect 14395 787 14473 833
rect 14519 787 14597 833
rect 14643 787 14721 833
rect 14767 787 15064 833
rect 14214 709 15064 787
rect 14214 663 14225 709
rect 14271 663 14349 709
rect 14395 663 14473 709
rect 14519 663 14597 709
rect 14643 663 14721 709
rect 14767 663 15064 709
rect 14214 496 15064 663
rect 0 338 122 496
rect 14942 338 15064 496
<< via1 >>
rect 2522 56786 2574 56790
rect 2646 56786 2698 56790
rect 2770 56786 2822 56790
rect 2894 56786 2946 56790
rect 3018 56786 3070 56790
rect 3142 56786 3194 56790
rect 3266 56786 3318 56790
rect 3390 56786 3442 56790
rect 3514 56786 3566 56790
rect 3638 56786 3690 56790
rect 3762 56786 3814 56790
rect 3886 56786 3938 56790
rect 4010 56786 4062 56790
rect 4134 56786 4186 56790
rect 4258 56786 4310 56790
rect 4382 56786 4434 56790
rect 4506 56786 4558 56790
rect 4630 56786 4682 56790
rect 4754 56786 4806 56790
rect 4878 56786 4930 56790
rect 5002 56786 5054 56790
rect 5126 56786 5178 56790
rect 5250 56786 5302 56790
rect 5374 56786 5426 56790
rect 5498 56786 5550 56790
rect 5622 56786 5674 56790
rect 5746 56786 5798 56790
rect 5870 56786 5922 56790
rect 5994 56786 6046 56790
rect 6118 56786 6170 56790
rect 6242 56786 6294 56790
rect 6366 56786 6418 56790
rect 6490 56786 6542 56790
rect 6614 56786 6666 56790
rect 6738 56786 6790 56790
rect 6862 56786 6914 56790
rect 6986 56786 7038 56790
rect 7110 56786 7162 56790
rect 7234 56786 7286 56790
rect 7358 56786 7410 56790
rect 7482 56786 7534 56790
rect 7606 56786 7658 56790
rect 7730 56786 7782 56790
rect 7854 56786 7906 56790
rect 7978 56786 8030 56790
rect 8102 56786 8154 56790
rect 8226 56786 8278 56790
rect 8350 56786 8402 56790
rect 8474 56786 8526 56790
rect 8598 56786 8650 56790
rect 8722 56786 8774 56790
rect 8846 56786 8898 56790
rect 8970 56786 9022 56790
rect 9094 56786 9146 56790
rect 9218 56786 9270 56790
rect 9342 56786 9394 56790
rect 9466 56786 9518 56790
rect 9590 56786 9642 56790
rect 9714 56786 9766 56790
rect 9838 56786 9890 56790
rect 9962 56786 10014 56790
rect 10086 56786 10138 56790
rect 10210 56786 10262 56790
rect 10334 56786 10386 56790
rect 10458 56786 10510 56790
rect 10582 56786 10634 56790
rect 10706 56786 10758 56790
rect 10830 56786 10882 56790
rect 10954 56786 11006 56790
rect 11078 56786 11130 56790
rect 11202 56786 11254 56790
rect 11326 56786 11378 56790
rect 11450 56786 11502 56790
rect 11574 56786 11626 56790
rect 11698 56786 11750 56790
rect 11822 56786 11874 56790
rect 11946 56786 11998 56790
rect 12070 56786 12122 56790
rect 12194 56786 12246 56790
rect 12318 56786 12370 56790
rect 12442 56786 12494 56790
rect 12566 56786 12618 56790
rect 12690 56786 12742 56790
rect 12814 56786 12866 56790
rect 12938 56786 12990 56790
rect 13062 56786 13114 56790
rect 13186 56786 13238 56790
rect 13310 56786 13362 56790
rect 13434 56786 13486 56790
rect 13558 56786 13610 56790
rect 2522 56738 2574 56786
rect 2646 56738 2698 56786
rect 2770 56738 2822 56786
rect 2894 56738 2946 56786
rect 3018 56738 3070 56786
rect 3142 56738 3194 56786
rect 3266 56738 3318 56786
rect 3390 56738 3442 56786
rect 3514 56738 3566 56786
rect 3638 56738 3690 56786
rect 3762 56738 3814 56786
rect 3886 56738 3938 56786
rect 4010 56738 4062 56786
rect 4134 56738 4186 56786
rect 4258 56738 4310 56786
rect 4382 56738 4434 56786
rect 4506 56738 4558 56786
rect 4630 56738 4682 56786
rect 4754 56738 4806 56786
rect 4878 56738 4930 56786
rect 5002 56738 5054 56786
rect 5126 56738 5178 56786
rect 5250 56738 5302 56786
rect 5374 56738 5426 56786
rect 5498 56738 5550 56786
rect 5622 56738 5674 56786
rect 5746 56738 5798 56786
rect 5870 56738 5922 56786
rect 5994 56738 6046 56786
rect 6118 56738 6170 56786
rect 6242 56738 6294 56786
rect 6366 56738 6418 56786
rect 6490 56738 6542 56786
rect 6614 56738 6666 56786
rect 6738 56738 6790 56786
rect 6862 56738 6914 56786
rect 6986 56738 7038 56786
rect 7110 56738 7162 56786
rect 7234 56738 7286 56786
rect 7358 56738 7410 56786
rect 7482 56738 7534 56786
rect 7606 56738 7658 56786
rect 7730 56738 7782 56786
rect 7854 56738 7906 56786
rect 7978 56738 8030 56786
rect 8102 56738 8154 56786
rect 8226 56738 8278 56786
rect 8350 56738 8402 56786
rect 8474 56738 8526 56786
rect 8598 56738 8650 56786
rect 8722 56738 8774 56786
rect 8846 56738 8898 56786
rect 8970 56738 9022 56786
rect 9094 56738 9146 56786
rect 9218 56738 9270 56786
rect 9342 56738 9394 56786
rect 9466 56738 9518 56786
rect 9590 56738 9642 56786
rect 9714 56738 9766 56786
rect 9838 56738 9890 56786
rect 9962 56738 10014 56786
rect 10086 56738 10138 56786
rect 10210 56738 10262 56786
rect 10334 56738 10386 56786
rect 10458 56738 10510 56786
rect 10582 56738 10634 56786
rect 10706 56738 10758 56786
rect 10830 56738 10882 56786
rect 10954 56738 11006 56786
rect 11078 56738 11130 56786
rect 11202 56738 11254 56786
rect 11326 56738 11378 56786
rect 11450 56738 11502 56786
rect 11574 56738 11626 56786
rect 11698 56738 11750 56786
rect 11822 56738 11874 56786
rect 11946 56738 11998 56786
rect 12070 56738 12122 56786
rect 12194 56738 12246 56786
rect 12318 56738 12370 56786
rect 12442 56738 12494 56786
rect 12566 56738 12618 56786
rect 12690 56738 12742 56786
rect 12814 56738 12866 56786
rect 12938 56738 12990 56786
rect 13062 56738 13114 56786
rect 13186 56738 13238 56786
rect 13310 56738 13362 56786
rect 13434 56738 13486 56786
rect 13558 56738 13610 56786
rect 2522 56614 2574 56666
rect 2646 56614 2698 56666
rect 2770 56614 2822 56666
rect 2894 56614 2946 56666
rect 3018 56614 3070 56666
rect 3142 56614 3194 56666
rect 3266 56614 3318 56666
rect 3390 56614 3442 56666
rect 3514 56614 3566 56666
rect 3638 56614 3690 56666
rect 3762 56614 3814 56666
rect 3886 56614 3938 56666
rect 4010 56614 4062 56666
rect 4134 56614 4186 56666
rect 4258 56614 4310 56666
rect 4382 56614 4434 56666
rect 4506 56614 4558 56666
rect 4630 56614 4682 56666
rect 4754 56614 4806 56666
rect 4878 56614 4930 56666
rect 5002 56614 5054 56666
rect 5126 56614 5178 56666
rect 5250 56614 5302 56666
rect 5374 56614 5426 56666
rect 5498 56614 5550 56666
rect 5622 56614 5674 56666
rect 5746 56614 5798 56666
rect 5870 56614 5922 56666
rect 5994 56614 6046 56666
rect 6118 56614 6170 56666
rect 6242 56614 6294 56666
rect 6366 56614 6418 56666
rect 6490 56614 6542 56666
rect 6614 56614 6666 56666
rect 6738 56614 6790 56666
rect 6862 56614 6914 56666
rect 6986 56614 7038 56666
rect 7110 56614 7162 56666
rect 7234 56614 7286 56666
rect 7358 56614 7410 56666
rect 7482 56614 7534 56666
rect 7606 56614 7658 56666
rect 7730 56614 7782 56666
rect 7854 56614 7906 56666
rect 7978 56614 8030 56666
rect 8102 56614 8154 56666
rect 8226 56614 8278 56666
rect 8350 56614 8402 56666
rect 8474 56614 8526 56666
rect 8598 56614 8650 56666
rect 8722 56614 8774 56666
rect 8846 56614 8898 56666
rect 8970 56614 9022 56666
rect 9094 56614 9146 56666
rect 9218 56614 9270 56666
rect 9342 56614 9394 56666
rect 9466 56614 9518 56666
rect 9590 56614 9642 56666
rect 9714 56614 9766 56666
rect 9838 56614 9890 56666
rect 9962 56614 10014 56666
rect 10086 56614 10138 56666
rect 10210 56614 10262 56666
rect 10334 56614 10386 56666
rect 10458 56614 10510 56666
rect 10582 56614 10634 56666
rect 10706 56614 10758 56666
rect 10830 56614 10882 56666
rect 10954 56614 11006 56666
rect 11078 56614 11130 56666
rect 11202 56614 11254 56666
rect 11326 56614 11378 56666
rect 11450 56614 11502 56666
rect 11574 56614 11626 56666
rect 11698 56614 11750 56666
rect 11822 56614 11874 56666
rect 11946 56614 11998 56666
rect 12070 56614 12122 56666
rect 12194 56614 12246 56666
rect 12318 56614 12370 56666
rect 12442 56614 12494 56666
rect 12566 56614 12618 56666
rect 12690 56614 12742 56666
rect 12814 56614 12866 56666
rect 12938 56614 12990 56666
rect 13062 56614 13114 56666
rect 13186 56614 13238 56666
rect 13310 56614 13362 56666
rect 13434 56614 13486 56666
rect 13558 56614 13610 56666
rect 2522 56490 2574 56542
rect 2646 56490 2698 56542
rect 2770 56494 2822 56542
rect 2894 56494 2946 56542
rect 3018 56494 3070 56542
rect 3142 56494 3194 56542
rect 3266 56494 3318 56542
rect 3390 56494 3442 56542
rect 3514 56494 3566 56542
rect 3638 56494 3690 56542
rect 2770 56490 2797 56494
rect 2797 56490 2822 56494
rect 2894 56490 2946 56494
rect 3018 56490 3070 56494
rect 3142 56490 3194 56494
rect 3266 56490 3318 56494
rect 3390 56490 3442 56494
rect 3514 56490 3566 56494
rect 3638 56490 3690 56494
rect 3762 56490 3814 56542
rect 3886 56490 3938 56542
rect 4010 56490 4062 56542
rect 4134 56490 4186 56542
rect 4258 56494 4310 56542
rect 4382 56494 4434 56542
rect 4506 56494 4558 56542
rect 4630 56494 4682 56542
rect 4754 56494 4806 56542
rect 4878 56494 4930 56542
rect 5002 56494 5054 56542
rect 5126 56494 5178 56542
rect 4258 56490 4297 56494
rect 4297 56490 4310 56494
rect 4382 56490 4434 56494
rect 4506 56490 4558 56494
rect 4630 56490 4682 56494
rect 4754 56490 4806 56494
rect 4878 56490 4930 56494
rect 5002 56490 5054 56494
rect 5126 56490 5178 56494
rect 5250 56490 5302 56542
rect 5374 56490 5426 56542
rect 5498 56490 5550 56542
rect 5622 56490 5674 56542
rect 5746 56494 5798 56542
rect 5870 56494 5922 56542
rect 5994 56494 6046 56542
rect 6118 56494 6170 56542
rect 6242 56494 6294 56542
rect 6366 56494 6418 56542
rect 6490 56494 6542 56542
rect 6614 56494 6666 56542
rect 5746 56490 5797 56494
rect 5797 56490 5798 56494
rect 5870 56490 5922 56494
rect 5994 56490 6046 56494
rect 6118 56490 6170 56494
rect 6242 56490 6294 56494
rect 6366 56490 6418 56494
rect 6490 56490 6542 56494
rect 6614 56490 6666 56494
rect 6738 56490 6790 56542
rect 6862 56490 6914 56542
rect 6986 56490 7038 56542
rect 7110 56490 7162 56542
rect 7234 56490 7286 56542
rect 7358 56494 7410 56542
rect 7482 56494 7534 56542
rect 7606 56494 7658 56542
rect 7730 56494 7782 56542
rect 7854 56494 7906 56542
rect 7978 56494 8030 56542
rect 8102 56494 8154 56542
rect 7358 56490 7410 56494
rect 7482 56490 7534 56494
rect 7606 56490 7658 56494
rect 7730 56490 7782 56494
rect 7854 56490 7906 56494
rect 7978 56490 8030 56494
rect 8102 56490 8154 56494
rect 8226 56490 8278 56542
rect 8350 56490 8402 56542
rect 8474 56490 8526 56542
rect 8598 56490 8650 56542
rect 8722 56490 8774 56542
rect 8846 56494 8898 56542
rect 8970 56494 9022 56542
rect 9094 56494 9146 56542
rect 9218 56494 9270 56542
rect 9342 56494 9394 56542
rect 9466 56494 9518 56542
rect 9590 56494 9642 56542
rect 9714 56494 9766 56542
rect 8846 56490 8898 56494
rect 8970 56490 9022 56494
rect 9094 56490 9146 56494
rect 9218 56490 9270 56494
rect 9342 56490 9394 56494
rect 9466 56490 9518 56494
rect 9590 56490 9642 56494
rect 9714 56490 9723 56494
rect 9723 56490 9766 56494
rect 9838 56490 9890 56542
rect 9962 56490 10014 56542
rect 10086 56490 10138 56542
rect 10210 56490 10262 56542
rect 10334 56494 10386 56542
rect 10458 56494 10510 56542
rect 10582 56494 10634 56542
rect 10706 56494 10758 56542
rect 10830 56494 10882 56542
rect 10954 56494 11006 56542
rect 11078 56494 11130 56542
rect 11202 56494 11254 56542
rect 10334 56490 10386 56494
rect 10458 56490 10510 56494
rect 10582 56490 10634 56494
rect 10706 56490 10758 56494
rect 10830 56490 10882 56494
rect 10954 56490 11006 56494
rect 11078 56490 11130 56494
rect 11202 56490 11223 56494
rect 11223 56490 11254 56494
rect 11326 56490 11378 56542
rect 11450 56490 11502 56542
rect 11574 56490 11626 56542
rect 11698 56490 11750 56542
rect 11822 56494 11874 56542
rect 11946 56494 11998 56542
rect 12070 56494 12122 56542
rect 12194 56494 12246 56542
rect 12318 56494 12370 56542
rect 12442 56494 12494 56542
rect 12566 56494 12618 56542
rect 12690 56494 12742 56542
rect 11822 56490 11874 56494
rect 11946 56490 11998 56494
rect 12070 56490 12122 56494
rect 12194 56490 12246 56494
rect 12318 56490 12370 56494
rect 12442 56490 12494 56494
rect 12566 56490 12618 56494
rect 12690 56490 12723 56494
rect 12723 56490 12742 56494
rect 12814 56490 12866 56542
rect 12938 56490 12990 56542
rect 13062 56490 13114 56542
rect 13186 56490 13238 56542
rect 13310 56494 13362 56542
rect 13434 56494 13486 56542
rect 13558 56494 13610 56542
rect 13310 56490 13362 56494
rect 13434 56490 13486 56494
rect 13558 56490 13610 56494
rect 2682 56320 2727 56345
rect 2727 56320 2838 56345
rect 2682 56218 2838 56320
rect 2682 56189 2727 56218
rect 2727 56189 2838 56218
rect 3682 56320 3793 56345
rect 3793 56320 3838 56345
rect 3682 56218 3838 56320
rect 3682 56189 3793 56218
rect 3793 56189 3838 56218
rect 4182 56320 4227 56345
rect 4227 56320 4338 56345
rect 4182 56218 4338 56320
rect 4182 56189 4227 56218
rect 4227 56189 4338 56218
rect 5182 56320 5293 56345
rect 5293 56320 5338 56345
rect 5182 56218 5338 56320
rect 5182 56189 5293 56218
rect 5293 56189 5338 56218
rect 5682 56320 5727 56345
rect 5727 56320 5838 56345
rect 5682 56218 5838 56320
rect 5682 56189 5727 56218
rect 5727 56189 5838 56218
rect 6682 56320 6793 56345
rect 6793 56320 6838 56345
rect 6682 56218 6838 56320
rect 6682 56189 6793 56218
rect 6793 56189 6838 56218
rect 7182 56320 7227 56345
rect 7227 56320 7338 56345
rect 7182 56218 7338 56320
rect 7182 56189 7227 56218
rect 7227 56189 7338 56218
rect 8182 56320 8293 56345
rect 8293 56320 8338 56345
rect 8182 56218 8338 56320
rect 8182 56189 8293 56218
rect 8293 56189 8338 56218
rect 8682 56320 8727 56345
rect 8727 56320 8838 56345
rect 8682 56218 8838 56320
rect 8682 56189 8727 56218
rect 8727 56189 8838 56218
rect 9682 56320 9793 56345
rect 9793 56320 9838 56345
rect 9682 56218 9838 56320
rect 9682 56189 9793 56218
rect 9793 56189 9838 56218
rect 10182 56320 10227 56345
rect 10227 56320 10338 56345
rect 10182 56218 10338 56320
rect 10182 56189 10227 56218
rect 10227 56189 10338 56218
rect 11182 56320 11293 56345
rect 11293 56320 11338 56345
rect 11182 56218 11338 56320
rect 11182 56189 11293 56218
rect 11293 56189 11338 56218
rect 11682 56320 11727 56345
rect 11727 56320 11838 56345
rect 11682 56218 11838 56320
rect 11682 56189 11727 56218
rect 11727 56189 11838 56218
rect 12682 56320 12793 56345
rect 12793 56320 12838 56345
rect 12682 56218 12838 56320
rect 12682 56189 12793 56218
rect 12793 56189 12838 56218
rect 13182 56320 13227 56345
rect 13227 56320 13338 56345
rect 13182 56218 13338 56320
rect 13182 56189 13227 56218
rect 13227 56189 13338 56218
rect 14392 56189 14548 56345
rect 2522 55996 2574 56048
rect 2646 55996 2698 56048
rect 2770 56044 2797 56048
rect 2797 56044 2822 56048
rect 2894 56044 2946 56048
rect 3018 56044 3070 56048
rect 3142 56044 3194 56048
rect 3266 56044 3318 56048
rect 3390 56044 3442 56048
rect 3514 56044 3566 56048
rect 3638 56044 3690 56048
rect 2770 55996 2822 56044
rect 2894 55996 2946 56044
rect 3018 55996 3070 56044
rect 3142 55996 3194 56044
rect 3266 55996 3318 56044
rect 3390 55996 3442 56044
rect 3514 55996 3566 56044
rect 3638 55996 3690 56044
rect 3762 55996 3814 56048
rect 3886 55996 3938 56048
rect 4010 55996 4062 56048
rect 4134 55996 4186 56048
rect 4258 56044 4297 56048
rect 4297 56044 4310 56048
rect 4382 56044 4434 56048
rect 4506 56044 4558 56048
rect 4630 56044 4682 56048
rect 4754 56044 4806 56048
rect 4878 56044 4930 56048
rect 5002 56044 5054 56048
rect 5126 56044 5178 56048
rect 4258 55996 4310 56044
rect 4382 55996 4434 56044
rect 4506 55996 4558 56044
rect 4630 55996 4682 56044
rect 4754 55996 4806 56044
rect 4878 55996 4930 56044
rect 5002 55996 5054 56044
rect 5126 55996 5178 56044
rect 5250 55996 5302 56048
rect 5374 55996 5426 56048
rect 5498 55996 5550 56048
rect 5622 55996 5674 56048
rect 5746 56044 5797 56048
rect 5797 56044 5798 56048
rect 5870 56044 5922 56048
rect 5994 56044 6046 56048
rect 6118 56044 6170 56048
rect 6242 56044 6294 56048
rect 6366 56044 6418 56048
rect 6490 56044 6542 56048
rect 6614 56044 6666 56048
rect 5746 55996 5798 56044
rect 5870 55996 5922 56044
rect 5994 55996 6046 56044
rect 6118 55996 6170 56044
rect 6242 55996 6294 56044
rect 6366 55996 6418 56044
rect 6490 55996 6542 56044
rect 6614 55996 6666 56044
rect 6738 55996 6790 56048
rect 6862 55996 6914 56048
rect 6986 55996 7038 56048
rect 7110 55996 7162 56048
rect 7234 55996 7286 56048
rect 7358 56044 7410 56048
rect 7482 56044 7534 56048
rect 7606 56044 7658 56048
rect 7730 56044 7782 56048
rect 7854 56044 7906 56048
rect 7978 56044 8030 56048
rect 8102 56044 8154 56048
rect 7358 55996 7410 56044
rect 7482 55996 7534 56044
rect 7606 55996 7658 56044
rect 7730 55996 7782 56044
rect 7854 55996 7906 56044
rect 7978 55996 8030 56044
rect 8102 55996 8154 56044
rect 8226 55996 8278 56048
rect 8350 55996 8402 56048
rect 8474 55996 8526 56048
rect 8598 55996 8650 56048
rect 8722 55996 8774 56048
rect 8846 56044 8898 56048
rect 8970 56044 9022 56048
rect 9094 56044 9146 56048
rect 9218 56044 9270 56048
rect 9342 56044 9394 56048
rect 9466 56044 9518 56048
rect 9590 56044 9642 56048
rect 9714 56044 9723 56048
rect 9723 56044 9766 56048
rect 8846 55996 8898 56044
rect 8970 55996 9022 56044
rect 9094 55996 9146 56044
rect 9218 55996 9270 56044
rect 9342 55996 9394 56044
rect 9466 55996 9518 56044
rect 9590 55996 9642 56044
rect 9714 55996 9766 56044
rect 9838 55996 9890 56048
rect 9962 55996 10014 56048
rect 10086 55996 10138 56048
rect 10210 55996 10262 56048
rect 10334 56044 10386 56048
rect 10458 56044 10510 56048
rect 10582 56044 10634 56048
rect 10706 56044 10758 56048
rect 10830 56044 10882 56048
rect 10954 56044 11006 56048
rect 11078 56044 11130 56048
rect 11202 56044 11223 56048
rect 11223 56044 11254 56048
rect 10334 55996 10386 56044
rect 10458 55996 10510 56044
rect 10582 55996 10634 56044
rect 10706 55996 10758 56044
rect 10830 55996 10882 56044
rect 10954 55996 11006 56044
rect 11078 55996 11130 56044
rect 11202 55996 11254 56044
rect 11326 55996 11378 56048
rect 11450 55996 11502 56048
rect 11574 55996 11626 56048
rect 11698 55996 11750 56048
rect 11822 56044 11874 56048
rect 11946 56044 11998 56048
rect 12070 56044 12122 56048
rect 12194 56044 12246 56048
rect 12318 56044 12370 56048
rect 12442 56044 12494 56048
rect 12566 56044 12618 56048
rect 12690 56044 12723 56048
rect 12723 56044 12742 56048
rect 11822 55996 11874 56044
rect 11946 55996 11998 56044
rect 12070 55996 12122 56044
rect 12194 55996 12246 56044
rect 12318 55996 12370 56044
rect 12442 55996 12494 56044
rect 12566 55996 12618 56044
rect 12690 55996 12742 56044
rect 12814 55996 12866 56048
rect 12938 55996 12990 56048
rect 13062 55996 13114 56048
rect 13186 55996 13238 56048
rect 13310 56044 13362 56048
rect 13434 56044 13486 56048
rect 13558 56044 13610 56048
rect 13310 55996 13362 56044
rect 13434 55996 13486 56044
rect 13558 55996 13610 56044
rect 2522 55872 2574 55924
rect 2646 55872 2698 55924
rect 2770 55872 2822 55924
rect 2894 55872 2946 55924
rect 3018 55872 3070 55924
rect 3142 55872 3194 55924
rect 3266 55872 3318 55924
rect 3390 55872 3442 55924
rect 3514 55872 3566 55924
rect 3638 55872 3690 55924
rect 3762 55872 3814 55924
rect 3886 55872 3938 55924
rect 4010 55872 4062 55924
rect 4134 55872 4186 55924
rect 4258 55872 4310 55924
rect 4382 55872 4434 55924
rect 4506 55872 4558 55924
rect 4630 55872 4682 55924
rect 4754 55872 4806 55924
rect 4878 55872 4930 55924
rect 5002 55872 5054 55924
rect 5126 55872 5178 55924
rect 5250 55872 5302 55924
rect 5374 55872 5426 55924
rect 5498 55872 5550 55924
rect 5622 55872 5674 55924
rect 5746 55872 5798 55924
rect 5870 55872 5922 55924
rect 5994 55872 6046 55924
rect 6118 55872 6170 55924
rect 6242 55872 6294 55924
rect 6366 55872 6418 55924
rect 6490 55872 6542 55924
rect 6614 55872 6666 55924
rect 6738 55872 6790 55924
rect 6862 55872 6914 55924
rect 6986 55872 7038 55924
rect 7110 55872 7162 55924
rect 7234 55872 7286 55924
rect 7358 55872 7410 55924
rect 7482 55872 7534 55924
rect 7606 55872 7658 55924
rect 7730 55872 7782 55924
rect 7854 55872 7906 55924
rect 7978 55872 8030 55924
rect 8102 55872 8154 55924
rect 8226 55872 8278 55924
rect 8350 55872 8402 55924
rect 8474 55872 8526 55924
rect 8598 55872 8650 55924
rect 8722 55872 8774 55924
rect 8846 55872 8898 55924
rect 8970 55872 9022 55924
rect 9094 55872 9146 55924
rect 9218 55872 9270 55924
rect 9342 55872 9394 55924
rect 9466 55872 9518 55924
rect 9590 55872 9642 55924
rect 9714 55872 9766 55924
rect 9838 55872 9890 55924
rect 9962 55872 10014 55924
rect 10086 55872 10138 55924
rect 10210 55872 10262 55924
rect 10334 55872 10386 55924
rect 10458 55872 10510 55924
rect 10582 55872 10634 55924
rect 10706 55872 10758 55924
rect 10830 55872 10882 55924
rect 10954 55872 11006 55924
rect 11078 55872 11130 55924
rect 11202 55872 11254 55924
rect 11326 55872 11378 55924
rect 11450 55872 11502 55924
rect 11574 55872 11626 55924
rect 11698 55872 11750 55924
rect 11822 55872 11874 55924
rect 11946 55872 11998 55924
rect 12070 55872 12122 55924
rect 12194 55872 12246 55924
rect 12318 55872 12370 55924
rect 12442 55872 12494 55924
rect 12566 55872 12618 55924
rect 12690 55872 12742 55924
rect 12814 55872 12866 55924
rect 12938 55872 12990 55924
rect 13062 55872 13114 55924
rect 13186 55872 13238 55924
rect 13310 55872 13362 55924
rect 13434 55872 13486 55924
rect 13558 55872 13610 55924
rect 1466 55374 1518 55530
rect 1608 55374 1660 55530
rect 2522 55752 2574 55800
rect 2646 55752 2698 55800
rect 2770 55752 2822 55800
rect 2894 55752 2946 55800
rect 3018 55752 3070 55800
rect 3142 55752 3194 55800
rect 3266 55752 3318 55800
rect 3390 55752 3442 55800
rect 3514 55752 3566 55800
rect 3638 55752 3690 55800
rect 3762 55752 3814 55800
rect 3886 55752 3938 55800
rect 4010 55752 4062 55800
rect 4134 55752 4186 55800
rect 4258 55752 4310 55800
rect 4382 55752 4434 55800
rect 4506 55752 4558 55800
rect 4630 55752 4682 55800
rect 4754 55752 4806 55800
rect 4878 55752 4930 55800
rect 5002 55752 5054 55800
rect 5126 55752 5178 55800
rect 5250 55752 5302 55800
rect 5374 55752 5426 55800
rect 5498 55752 5550 55800
rect 5622 55752 5674 55800
rect 5746 55752 5798 55800
rect 5870 55752 5922 55800
rect 5994 55752 6046 55800
rect 6118 55752 6170 55800
rect 6242 55752 6294 55800
rect 6366 55752 6418 55800
rect 6490 55752 6542 55800
rect 6614 55752 6666 55800
rect 6738 55752 6790 55800
rect 6862 55752 6914 55800
rect 6986 55752 7038 55800
rect 7110 55752 7162 55800
rect 7234 55752 7286 55800
rect 7358 55752 7410 55800
rect 7482 55752 7534 55800
rect 7606 55752 7658 55800
rect 7730 55752 7782 55800
rect 7854 55752 7906 55800
rect 7978 55752 8030 55800
rect 8102 55752 8154 55800
rect 8226 55752 8278 55800
rect 8350 55752 8402 55800
rect 8474 55752 8526 55800
rect 8598 55752 8650 55800
rect 8722 55752 8774 55800
rect 8846 55752 8898 55800
rect 8970 55752 9022 55800
rect 9094 55752 9146 55800
rect 9218 55752 9270 55800
rect 9342 55752 9394 55800
rect 9466 55752 9518 55800
rect 9590 55752 9642 55800
rect 9714 55752 9766 55800
rect 9838 55752 9890 55800
rect 9962 55752 10014 55800
rect 10086 55752 10138 55800
rect 10210 55752 10262 55800
rect 10334 55752 10386 55800
rect 10458 55752 10510 55800
rect 10582 55752 10634 55800
rect 10706 55752 10758 55800
rect 10830 55752 10882 55800
rect 10954 55752 11006 55800
rect 11078 55752 11130 55800
rect 11202 55752 11254 55800
rect 11326 55752 11378 55800
rect 11450 55752 11502 55800
rect 11574 55752 11626 55800
rect 11698 55752 11750 55800
rect 11822 55752 11874 55800
rect 11946 55752 11998 55800
rect 12070 55752 12122 55800
rect 12194 55752 12246 55800
rect 12318 55752 12370 55800
rect 12442 55752 12494 55800
rect 12566 55752 12618 55800
rect 12690 55752 12742 55800
rect 12814 55752 12866 55800
rect 12938 55752 12990 55800
rect 13062 55752 13114 55800
rect 13186 55752 13238 55800
rect 13310 55752 13362 55800
rect 13434 55752 13486 55800
rect 13558 55752 13610 55800
rect 2522 55748 2574 55752
rect 2646 55748 2698 55752
rect 2770 55748 2822 55752
rect 2894 55748 2946 55752
rect 3018 55748 3070 55752
rect 3142 55748 3194 55752
rect 3266 55748 3318 55752
rect 3390 55748 3442 55752
rect 3514 55748 3566 55752
rect 3638 55748 3690 55752
rect 3762 55748 3814 55752
rect 3886 55748 3938 55752
rect 4010 55748 4062 55752
rect 4134 55748 4186 55752
rect 4258 55748 4310 55752
rect 4382 55748 4434 55752
rect 4506 55748 4558 55752
rect 4630 55748 4682 55752
rect 4754 55748 4806 55752
rect 4878 55748 4930 55752
rect 5002 55748 5054 55752
rect 5126 55748 5178 55752
rect 5250 55748 5302 55752
rect 5374 55748 5426 55752
rect 5498 55748 5550 55752
rect 5622 55748 5674 55752
rect 5746 55748 5798 55752
rect 5870 55748 5922 55752
rect 5994 55748 6046 55752
rect 6118 55748 6170 55752
rect 6242 55748 6294 55752
rect 6366 55748 6418 55752
rect 6490 55748 6542 55752
rect 6614 55748 6666 55752
rect 6738 55748 6790 55752
rect 6862 55748 6914 55752
rect 6986 55748 7038 55752
rect 7110 55748 7162 55752
rect 7234 55748 7286 55752
rect 7358 55748 7410 55752
rect 7482 55748 7534 55752
rect 7606 55748 7658 55752
rect 7730 55748 7782 55752
rect 7854 55748 7906 55752
rect 7978 55748 8030 55752
rect 8102 55748 8154 55752
rect 8226 55748 8278 55752
rect 8350 55748 8402 55752
rect 8474 55748 8526 55752
rect 8598 55748 8650 55752
rect 8722 55748 8774 55752
rect 8846 55748 8898 55752
rect 8970 55748 9022 55752
rect 9094 55748 9146 55752
rect 9218 55748 9270 55752
rect 9342 55748 9394 55752
rect 9466 55748 9518 55752
rect 9590 55748 9642 55752
rect 9714 55748 9766 55752
rect 9838 55748 9890 55752
rect 9962 55748 10014 55752
rect 10086 55748 10138 55752
rect 10210 55748 10262 55752
rect 10334 55748 10386 55752
rect 10458 55748 10510 55752
rect 10582 55748 10634 55752
rect 10706 55748 10758 55752
rect 10830 55748 10882 55752
rect 10954 55748 11006 55752
rect 11078 55748 11130 55752
rect 11202 55748 11254 55752
rect 11326 55748 11378 55752
rect 11450 55748 11502 55752
rect 11574 55748 11626 55752
rect 11698 55748 11750 55752
rect 11822 55748 11874 55752
rect 11946 55748 11998 55752
rect 12070 55748 12122 55752
rect 12194 55748 12246 55752
rect 12318 55748 12370 55752
rect 12442 55748 12494 55752
rect 12566 55748 12618 55752
rect 12690 55748 12742 55752
rect 12814 55748 12866 55752
rect 12938 55748 12990 55752
rect 13062 55748 13114 55752
rect 13186 55748 13238 55752
rect 13310 55748 13362 55752
rect 13434 55748 13486 55752
rect 13558 55748 13610 55752
rect 234 54673 286 54725
rect 358 54673 410 54725
rect 482 54673 534 54725
rect 234 54549 286 54601
rect 358 54549 410 54601
rect 482 54549 534 54601
rect 234 54425 286 54477
rect 358 54425 410 54477
rect 482 54425 534 54477
rect 3482 54471 3534 55459
rect 3705 54471 3757 55459
rect 4174 54471 4226 55459
rect 4770 54624 4822 55404
rect 4950 54624 5002 55404
rect 5438 54624 5490 55404
rect 5926 54624 5978 55404
rect 6108 54475 6160 55359
rect 6290 54624 6342 55404
rect 6778 54624 6830 55404
rect 7266 54624 7318 55404
rect 7446 54624 7498 55404
rect 8042 54471 8094 55459
rect 8511 54471 8563 55459
rect 8726 54471 8778 55459
rect 8949 54471 9001 55459
rect 9418 54471 9470 55459
rect 10014 54624 10066 55404
rect 10194 54624 10246 55404
rect 10682 54624 10734 55404
rect 11170 54624 11222 55404
rect 11352 54475 11404 55359
rect 11534 54624 11586 55404
rect 12022 54624 12074 55404
rect 12510 54624 12562 55404
rect 12690 54624 12742 55404
rect 13286 54471 13338 55459
rect 234 53773 286 53825
rect 358 53773 410 53825
rect 482 53773 534 53825
rect 234 53649 286 53701
rect 358 53649 410 53701
rect 482 53649 534 53701
rect 234 53525 286 53577
rect 358 53525 410 53577
rect 482 53525 534 53577
rect 3482 53013 3534 54001
rect 4174 53013 4226 53793
rect 4770 53060 4822 53632
rect 4950 53060 5002 53632
rect 5438 53060 5490 53632
rect 5926 53060 5978 53632
rect 6108 53013 6160 53897
rect 6290 53060 6342 53632
rect 6778 53060 6830 53632
rect 7266 53060 7318 53632
rect 7446 53060 7498 53632
rect 8042 53013 8094 53793
rect 8730 53013 8782 54001
rect 10014 53060 10066 53632
rect 10194 53060 10246 53632
rect 10682 53060 10734 53632
rect 11170 53060 11222 53632
rect 11352 53013 11404 53897
rect 11534 53060 11586 53632
rect 12022 53060 12074 53632
rect 12510 53060 12562 53632
rect 12690 53060 12742 53632
rect 13286 53013 13338 53793
rect 722 52585 1086 52637
rect 3378 52585 3534 52637
rect 3727 52585 3883 52637
rect 6450 52257 6918 52309
rect 7266 52257 7422 52309
rect 58 50880 110 52180
rect 14954 50880 15006 52180
rect 2540 49847 6128 49899
rect 7732 49847 8096 49899
rect 8434 49847 8798 49899
rect 3990 48864 4042 48916
rect 4114 48864 4166 48916
rect 4238 48864 4290 48916
rect 3990 48740 4042 48792
rect 4114 48740 4166 48792
rect 4238 48740 4290 48792
rect 3990 48616 4042 48668
rect 4114 48616 4166 48668
rect 4238 48616 4290 48668
rect 3990 48492 4042 48544
rect 4114 48492 4166 48544
rect 4238 48492 4290 48544
rect 3990 48368 4042 48420
rect 4114 48368 4166 48420
rect 4238 48368 4290 48420
rect 3990 48244 4042 48296
rect 4114 48244 4166 48296
rect 4238 48244 4290 48296
rect 3990 48120 4042 48172
rect 4114 48120 4166 48172
rect 4238 48120 4290 48172
rect 3990 47996 4042 48048
rect 4114 47996 4166 48048
rect 4238 47996 4290 48048
rect 3990 47872 4042 47924
rect 4114 47872 4166 47924
rect 4238 47872 4290 47924
rect 3990 47748 4042 47800
rect 4114 47748 4166 47800
rect 4238 47748 4290 47800
rect 3620 46326 3672 47418
rect 3197 45666 3353 46134
rect 4644 49002 4696 49054
rect 4768 49002 4820 49054
rect 4892 49002 4944 49054
rect 4644 48878 4696 48930
rect 4768 48878 4820 48930
rect 4892 48878 4944 48930
rect 4644 48754 4696 48806
rect 4768 48754 4820 48806
rect 4892 48754 4944 48806
rect 5531 48768 5895 49028
rect 7732 48768 8096 49028
rect 8434 48768 8798 49028
rect 4644 48630 4696 48682
rect 4768 48630 4820 48682
rect 4892 48630 4944 48682
rect 4644 48506 4696 48558
rect 4768 48506 4820 48558
rect 4892 48506 4944 48558
rect 4644 48382 4696 48434
rect 4768 48382 4820 48434
rect 4892 48382 4944 48434
rect 4644 48258 4696 48310
rect 4768 48258 4820 48310
rect 4892 48258 4944 48310
rect 4644 48134 4696 48186
rect 4768 48134 4820 48186
rect 4892 48134 4944 48186
rect 4644 48010 4696 48062
rect 4768 48010 4820 48062
rect 4892 48010 4944 48062
rect 10794 48002 10846 48990
rect 4644 47886 4696 47938
rect 4768 47886 4820 47938
rect 4892 47886 4944 47938
rect 4644 47762 4696 47814
rect 4768 47762 4820 47814
rect 4892 47762 4944 47814
rect 4644 47638 4696 47690
rect 4768 47638 4820 47690
rect 4892 47638 4944 47690
rect 4644 47514 4696 47566
rect 4768 47514 4820 47566
rect 4892 47514 4944 47566
rect 11608 47452 11660 47608
rect 11013 46624 11065 47404
rect 3981 45287 4033 45339
rect 4105 45287 4157 45339
rect 4229 45287 4281 45339
rect 3981 45163 4033 45215
rect 4105 45163 4157 45215
rect 4229 45163 4281 45215
rect 3981 45039 4033 45091
rect 4105 45039 4157 45091
rect 4229 45039 4281 45091
rect 3981 44915 4033 44967
rect 4105 44915 4157 44967
rect 4229 44915 4281 44967
rect 3981 44791 4033 44843
rect 4105 44791 4157 44843
rect 4229 44791 4281 44843
rect 3981 44667 4033 44719
rect 4105 44667 4157 44719
rect 4229 44667 4281 44719
rect 3981 44543 4033 44595
rect 4105 44543 4157 44595
rect 4229 44543 4281 44595
rect 3620 42880 3672 44180
rect 12437 43631 12593 43683
rect 3620 41280 3672 42580
rect 11517 41288 11569 41444
rect 1848 40648 3668 40700
rect 11149 40637 11201 40793
rect 11532 40815 11584 40971
rect 13108 42469 13160 42498
rect 13108 42423 13115 42469
rect 13115 42423 13160 42469
rect 13108 42357 13160 42423
rect 13108 42342 13115 42357
rect 13115 42342 13160 42357
rect 13544 42469 13596 42498
rect 13544 42423 13589 42469
rect 13589 42423 13596 42469
rect 13544 42357 13596 42423
rect 13544 42342 13589 42357
rect 13589 42342 13596 42357
rect 13108 41567 13115 41571
rect 13115 41567 13160 41571
rect 13108 41501 13160 41567
rect 13108 41455 13115 41501
rect 13115 41455 13160 41501
rect 13108 41415 13160 41455
rect 13544 41567 13589 41571
rect 13589 41567 13596 41571
rect 13544 41501 13596 41567
rect 13544 41455 13589 41501
rect 13589 41455 13596 41501
rect 13544 41415 13596 41455
rect 1925 40312 2081 40364
rect 4849 40312 5005 40364
rect 7065 40312 7221 40364
rect 10796 40312 10952 40364
rect 14070 40312 14122 40468
rect 1608 40176 1764 40228
rect 5578 40176 5734 40228
rect 11428 40176 11584 40228
rect 13674 40176 13830 40228
rect 10656 40040 10812 40092
rect 11996 40040 12152 40092
rect 13820 40040 13976 40092
rect 202 39884 566 39936
rect 2445 39892 4473 39944
rect 7900 39892 9720 39944
rect 12784 39892 13772 39944
rect 1783 38846 1835 39418
rect 5095 38846 5147 39418
rect 6061 38430 6113 39418
rect 7027 38846 7079 39418
rect 10339 38430 10391 39418
rect 10656 38520 10708 38676
rect 10900 38520 10952 38676
rect 11212 38430 11264 39418
rect 8305 38162 8357 38318
rect 58 36480 110 37780
rect 817 37154 869 38142
rect 2719 37413 2771 37569
rect 3207 37413 3259 37569
rect 3439 37154 3491 38142
rect 11532 38159 11584 38315
rect 3671 37413 3723 37569
rect 4159 37413 4211 37569
rect 6061 37154 6113 38142
rect 13315 38151 13367 38307
rect 8451 37413 8503 37569
rect 8683 37154 8735 38142
rect 8907 37413 8959 37569
rect 13451 37497 13503 37653
rect 10343 37146 11539 37198
rect 8451 36476 8503 36632
rect 13074 36476 13230 36528
rect 8305 36340 8461 36392
rect 12934 36340 13090 36392
rect 2088 36204 2452 36256
rect 4473 36204 4629 36256
rect 5822 36204 5978 36256
rect 8982 36204 9138 36256
rect 1834 36068 1990 36120
rect 3103 36068 3259 36120
rect 3671 36068 3827 36120
rect 6066 36068 6222 36120
rect 8842 36068 8998 36120
rect 2494 35932 2650 35984
rect 5406 35932 5562 35984
rect 9502 35932 9658 35984
rect 12518 35932 12674 35984
rect 1322 35796 1478 35848
rect 6578 35796 6734 35848
rect 8330 35796 8486 35848
rect 13586 35796 13742 35848
rect 3398 35660 3554 35712
rect 4502 35660 4658 35712
rect 10406 35660 10562 35712
rect 11510 35660 11666 35712
rect 13347 35660 13503 35712
rect 498 33756 550 35576
rect 736 34172 788 35576
rect 3104 34172 3156 35576
rect 1834 33909 1886 34065
rect 2078 33909 2130 34065
rect 2494 33909 2546 34065
rect 498 29685 550 33481
rect 4002 32924 4054 35576
rect 4900 34172 4952 35576
rect 8579 35524 8735 35576
rect 10112 34172 10164 35576
rect 5510 33909 5562 34065
rect 5926 33909 5978 34065
rect 6170 33909 6222 34065
rect 8842 33909 8894 34065
rect 9086 33909 9138 34065
rect 9502 33909 9554 34065
rect 11010 32924 11062 35576
rect 11908 34172 11960 35576
rect 14954 36480 15006 37780
rect 12518 33909 12570 34065
rect 12934 33909 12986 34065
rect 13178 33909 13230 34065
rect 980 30084 1032 32320
rect 1468 29944 1520 30308
rect 1712 29944 1764 30308
rect 2372 30084 2424 32320
rect 2788 30084 2840 32320
rect 3276 30708 3328 32320
rect 3764 30658 3816 32270
rect 4002 30635 4054 32455
rect 4240 30658 4292 32270
rect 4728 30708 4780 32320
rect 5216 30708 5268 32320
rect 5632 30708 5684 32320
rect 3032 30124 3084 30488
rect 3520 29944 3572 30308
rect 4484 30124 4536 30488
rect 4972 29944 5024 30308
rect 6536 29944 6588 30308
rect 6780 29944 6832 30308
rect 7024 30084 7076 32320
rect 7988 30084 8040 32320
rect 9380 30708 9432 32320
rect 9796 30708 9848 32320
rect 10284 30708 10336 32320
rect 10772 30658 10824 32270
rect 11010 30635 11062 32455
rect 11248 30658 11300 32270
rect 11736 30708 11788 32320
rect 8476 29944 8528 30308
rect 8720 29944 8772 30308
rect 10040 29944 10092 30308
rect 10528 30124 10580 30488
rect 11492 29944 11544 30308
rect 11980 30124 12032 30488
rect 12224 30084 12276 32320
rect 12640 30084 12692 32320
rect 13544 29944 13596 30308
rect 13788 29944 13840 30308
rect 14032 30084 14084 32320
rect 2012 29685 3312 29737
rect 11949 29685 13249 29737
rect 14514 29685 14566 33481
rect 1379 29395 1535 29447
rect 6444 29395 6600 29447
rect 8708 29395 8864 29447
rect 13531 29395 13687 29447
rect 1559 29215 1715 29267
rect 6688 29215 6844 29267
rect 8464 29215 8620 29267
rect 13351 29215 13507 29267
rect 3508 29008 3664 29060
rect 4167 28943 4219 29099
rect 4972 28943 5024 29099
rect 5926 28943 5978 29099
rect 9088 28943 9140 29099
rect 10042 28943 10094 29099
rect 10847 28943 10899 29099
rect 11402 29008 11558 29060
<< metal2 >>
rect 704 55060 780 57230
rect 1225 55060 1301 57230
rect 1886 56865 1962 56875
rect 1886 56809 1896 56865
rect 1952 56809 1962 56865
rect 1886 56723 1962 56809
rect 1886 56667 1896 56723
rect 1952 56667 1962 56723
rect 1886 56581 1962 56667
rect 1886 56525 1896 56581
rect 1952 56525 1962 56581
rect 1886 56439 1962 56525
rect 1886 56383 1896 56439
rect 1952 56383 1962 56439
rect 1886 56297 1962 56383
rect 1886 56241 1896 56297
rect 1952 56241 1962 56297
rect 1886 56155 1962 56241
rect 1886 56099 1896 56155
rect 1952 56099 1962 56155
rect 1886 56013 1962 56099
rect 1886 55957 1896 56013
rect 1952 55957 1962 56013
rect 1886 55871 1962 55957
rect 1886 55815 1896 55871
rect 1952 55815 1962 55871
rect 1886 55729 1962 55815
rect 1886 55673 1896 55729
rect 1952 55673 1962 55729
rect 1454 55530 1530 55542
rect 1454 55374 1466 55530
rect 1518 55374 1530 55530
rect 184 54725 584 54799
rect 184 54673 234 54725
rect 286 54673 358 54725
rect 410 54673 482 54725
rect 534 54673 584 54725
rect 184 54601 584 54673
rect 184 54549 234 54601
rect 286 54549 358 54601
rect 410 54549 482 54601
rect 534 54549 584 54601
rect 184 54477 584 54549
rect 184 54425 234 54477
rect 286 54425 358 54477
rect 410 54425 482 54477
rect 534 54425 584 54477
rect 184 53825 584 54425
rect 184 53773 234 53825
rect 286 53773 358 53825
rect 410 53773 482 53825
rect 534 53773 584 53825
rect 184 53701 584 53773
rect 184 53649 234 53701
rect 286 53649 358 53701
rect 410 53649 482 53701
rect 534 53649 584 53701
rect 184 53577 584 53649
rect 184 53525 234 53577
rect 286 53525 358 53577
rect 410 53525 482 53577
rect 534 53525 584 53577
rect 32 52197 122 52230
rect 32 52141 56 52197
rect 112 52141 122 52197
rect 32 52055 58 52141
rect 110 52055 122 52141
rect 32 51999 56 52055
rect 112 51999 122 52055
rect 32 51913 58 51999
rect 110 51913 122 51999
rect 32 51857 56 51913
rect 112 51857 122 51913
rect 32 51771 58 51857
rect 110 51771 122 51857
rect 32 51715 56 51771
rect 112 51715 122 51771
rect 32 51629 58 51715
rect 110 51629 122 51715
rect 32 51573 56 51629
rect 112 51573 122 51629
rect 32 51487 58 51573
rect 110 51487 122 51573
rect 32 51431 56 51487
rect 112 51431 122 51487
rect 32 51345 58 51431
rect 110 51345 122 51431
rect 32 51289 56 51345
rect 112 51289 122 51345
rect 32 51203 58 51289
rect 110 51203 122 51289
rect 32 51147 56 51203
rect 112 51147 122 51203
rect 32 51061 58 51147
rect 110 51061 122 51147
rect 32 51005 56 51061
rect 112 51005 122 51061
rect 32 50919 58 51005
rect 110 50919 122 51005
rect 32 50863 56 50919
rect 112 50863 122 50919
rect 32 50830 122 50863
rect 184 50597 584 53525
rect 184 50541 214 50597
rect 270 50541 356 50597
rect 412 50541 498 50597
rect 554 50541 584 50597
rect 184 50455 584 50541
rect 184 50399 214 50455
rect 270 50399 356 50455
rect 412 50399 498 50455
rect 554 50399 584 50455
rect 184 50313 584 50399
rect 184 50257 214 50313
rect 270 50257 356 50313
rect 412 50257 498 50313
rect 554 50257 584 50313
rect 184 50171 584 50257
rect 184 50115 214 50171
rect 270 50115 356 50171
rect 412 50115 498 50171
rect 554 50115 584 50171
rect 184 50029 584 50115
rect 184 49973 214 50029
rect 270 49973 356 50029
rect 412 49973 498 50029
rect 554 49973 584 50029
rect 184 49887 584 49973
rect 184 49831 214 49887
rect 270 49831 356 49887
rect 412 49831 498 49887
rect 554 49831 584 49887
rect 184 49745 584 49831
rect 184 49689 214 49745
rect 270 49689 356 49745
rect 412 49689 498 49745
rect 554 49689 584 49745
rect 184 49603 584 49689
rect 184 49547 214 49603
rect 270 49547 356 49603
rect 412 49547 498 49603
rect 554 49547 584 49603
rect 184 49461 584 49547
rect 184 49405 214 49461
rect 270 49405 356 49461
rect 412 49405 498 49461
rect 554 49405 584 49461
rect 184 49319 584 49405
rect 184 49263 214 49319
rect 270 49263 356 49319
rect 412 49263 498 49319
rect 554 49263 584 49319
rect 184 39936 584 49263
rect 184 39884 202 39936
rect 566 39884 584 39936
rect 184 39397 584 39884
rect 184 39341 214 39397
rect 270 39341 356 39397
rect 412 39341 498 39397
rect 554 39341 584 39397
rect 184 39255 584 39341
rect 184 39199 214 39255
rect 270 39199 356 39255
rect 412 39199 498 39255
rect 554 39199 584 39255
rect 184 39113 584 39199
rect 184 39057 214 39113
rect 270 39057 356 39113
rect 412 39057 498 39113
rect 554 39057 584 39113
rect 184 38971 584 39057
rect 184 38915 214 38971
rect 270 38915 356 38971
rect 412 38915 498 38971
rect 554 38915 584 38971
rect 184 38829 584 38915
rect 184 38773 214 38829
rect 270 38773 356 38829
rect 412 38773 498 38829
rect 554 38773 584 38829
rect 184 38687 584 38773
rect 184 38631 214 38687
rect 270 38631 356 38687
rect 412 38631 498 38687
rect 554 38631 584 38687
rect 184 38545 584 38631
rect 184 38489 214 38545
rect 270 38489 356 38545
rect 412 38489 498 38545
rect 554 38489 584 38545
rect 184 38403 584 38489
rect 184 38347 214 38403
rect 270 38347 356 38403
rect 412 38347 498 38403
rect 554 38347 584 38403
rect 184 38261 584 38347
rect 184 38205 214 38261
rect 270 38205 356 38261
rect 412 38205 498 38261
rect 554 38205 584 38261
rect 184 38119 584 38205
rect 184 38063 214 38119
rect 270 38063 356 38119
rect 412 38063 498 38119
rect 554 38063 584 38119
rect 184 38030 584 38063
rect 704 52637 1104 52649
rect 704 52585 722 52637
rect 1086 52585 1104 52637
rect 704 52197 1104 52585
rect 704 52141 734 52197
rect 790 52141 876 52197
rect 932 52141 1018 52197
rect 1074 52141 1104 52197
rect 704 52055 1104 52141
rect 704 51999 734 52055
rect 790 51999 876 52055
rect 932 51999 1018 52055
rect 1074 51999 1104 52055
rect 704 51913 1104 51999
rect 704 51857 734 51913
rect 790 51857 876 51913
rect 932 51857 1018 51913
rect 1074 51857 1104 51913
rect 704 51771 1104 51857
rect 704 51715 734 51771
rect 790 51715 876 51771
rect 932 51715 1018 51771
rect 1074 51715 1104 51771
rect 704 51629 1104 51715
rect 704 51573 734 51629
rect 790 51573 876 51629
rect 932 51573 1018 51629
rect 1074 51573 1104 51629
rect 704 51487 1104 51573
rect 704 51431 734 51487
rect 790 51431 876 51487
rect 932 51431 1018 51487
rect 1074 51431 1104 51487
rect 704 51345 1104 51431
rect 704 51289 734 51345
rect 790 51289 876 51345
rect 932 51289 1018 51345
rect 1074 51289 1104 51345
rect 704 51203 1104 51289
rect 704 51147 734 51203
rect 790 51147 876 51203
rect 932 51147 1018 51203
rect 1074 51147 1104 51203
rect 704 51061 1104 51147
rect 704 51005 734 51061
rect 790 51005 876 51061
rect 932 51005 1018 51061
rect 1074 51005 1104 51061
rect 704 50919 1104 51005
rect 704 50863 734 50919
rect 790 50863 876 50919
rect 932 50863 1018 50919
rect 1074 50863 1104 50919
rect 704 38142 1104 50863
rect 1454 40239 1530 55374
rect 1184 40163 1530 40239
rect 1596 55530 1672 55542
rect 1596 55374 1608 55530
rect 1660 55374 1672 55530
rect 1596 40240 1672 55374
rect 1886 53797 1962 55673
rect 1886 53741 1896 53797
rect 1952 53741 1962 53797
rect 1886 53655 1962 53741
rect 1886 53599 1896 53655
rect 1952 53599 1962 53655
rect 1886 53513 1962 53599
rect 1886 53457 1896 53513
rect 1952 53457 1962 53513
rect 1886 53371 1962 53457
rect 1886 53315 1896 53371
rect 1952 53315 1962 53371
rect 1886 53229 1962 53315
rect 1886 53173 1896 53229
rect 1952 53173 1962 53229
rect 2098 53296 2174 57230
rect 2309 54120 2385 57230
rect 2490 56810 13642 56820
rect 2490 56754 2500 56810
rect 2556 56790 2642 56810
rect 2698 56790 2784 56810
rect 2840 56790 2926 56810
rect 2982 56790 3068 56810
rect 3124 56790 3210 56810
rect 2574 56754 2642 56790
rect 2490 56738 2522 56754
rect 2574 56738 2646 56754
rect 2698 56738 2770 56790
rect 2840 56754 2894 56790
rect 2982 56754 3018 56790
rect 3124 56754 3142 56790
rect 2822 56738 2894 56754
rect 2946 56738 3018 56754
rect 3070 56738 3142 56754
rect 3194 56754 3210 56790
rect 3266 56790 3352 56810
rect 3408 56790 3494 56810
rect 3550 56790 3636 56810
rect 3692 56790 3778 56810
rect 3834 56790 3920 56810
rect 3976 56790 4062 56810
rect 3194 56738 3266 56754
rect 3318 56754 3352 56790
rect 3442 56754 3494 56790
rect 3566 56754 3636 56790
rect 3692 56754 3762 56790
rect 3834 56754 3886 56790
rect 3976 56754 4010 56790
rect 3318 56738 3390 56754
rect 3442 56738 3514 56754
rect 3566 56738 3638 56754
rect 3690 56738 3762 56754
rect 3814 56738 3886 56754
rect 3938 56738 4010 56754
rect 4118 56790 4204 56810
rect 4260 56790 4346 56810
rect 4402 56790 4488 56810
rect 4544 56790 4630 56810
rect 4686 56790 4772 56810
rect 4828 56790 4914 56810
rect 4970 56790 5056 56810
rect 4118 56754 4134 56790
rect 4062 56738 4134 56754
rect 4186 56754 4204 56790
rect 4310 56754 4346 56790
rect 4434 56754 4488 56790
rect 4186 56738 4258 56754
rect 4310 56738 4382 56754
rect 4434 56738 4506 56754
rect 4558 56738 4630 56790
rect 4686 56754 4754 56790
rect 4828 56754 4878 56790
rect 4970 56754 5002 56790
rect 4682 56738 4754 56754
rect 4806 56738 4878 56754
rect 4930 56738 5002 56754
rect 5054 56754 5056 56790
rect 5112 56790 5198 56810
rect 5254 56790 5340 56810
rect 5396 56790 5482 56810
rect 5538 56790 5624 56810
rect 5680 56790 5766 56810
rect 5822 56790 5908 56810
rect 5964 56790 6050 56810
rect 5112 56754 5126 56790
rect 5054 56738 5126 56754
rect 5178 56754 5198 56790
rect 5302 56754 5340 56790
rect 5426 56754 5482 56790
rect 5178 56738 5250 56754
rect 5302 56738 5374 56754
rect 5426 56738 5498 56754
rect 5550 56738 5622 56790
rect 5680 56754 5746 56790
rect 5822 56754 5870 56790
rect 5964 56754 5994 56790
rect 5674 56738 5746 56754
rect 5798 56738 5870 56754
rect 5922 56738 5994 56754
rect 6046 56754 6050 56790
rect 6106 56790 6192 56810
rect 6248 56790 6334 56810
rect 6390 56790 6476 56810
rect 6532 56790 6618 56810
rect 6674 56790 6760 56810
rect 6816 56790 6902 56810
rect 6958 56790 7044 56810
rect 6106 56754 6118 56790
rect 6046 56738 6118 56754
rect 6170 56754 6192 56790
rect 6294 56754 6334 56790
rect 6418 56754 6476 56790
rect 6170 56738 6242 56754
rect 6294 56738 6366 56754
rect 6418 56738 6490 56754
rect 6542 56738 6614 56790
rect 6674 56754 6738 56790
rect 6816 56754 6862 56790
rect 6958 56754 6986 56790
rect 6666 56738 6738 56754
rect 6790 56738 6862 56754
rect 6914 56738 6986 56754
rect 7038 56754 7044 56790
rect 7100 56790 7186 56810
rect 7242 56790 7328 56810
rect 7384 56790 7470 56810
rect 7526 56790 7612 56810
rect 7668 56790 7754 56810
rect 7810 56790 7896 56810
rect 7952 56790 8038 56810
rect 7100 56754 7110 56790
rect 7038 56738 7110 56754
rect 7162 56754 7186 56790
rect 7286 56754 7328 56790
rect 7410 56754 7470 56790
rect 7162 56738 7234 56754
rect 7286 56738 7358 56754
rect 7410 56738 7482 56754
rect 7534 56738 7606 56790
rect 7668 56754 7730 56790
rect 7810 56754 7854 56790
rect 7952 56754 7978 56790
rect 7658 56738 7730 56754
rect 7782 56738 7854 56754
rect 7906 56738 7978 56754
rect 8030 56754 8038 56790
rect 8094 56790 8180 56810
rect 8236 56790 8322 56810
rect 8378 56790 8464 56810
rect 8520 56790 8606 56810
rect 8662 56790 8748 56810
rect 8804 56790 8890 56810
rect 8946 56790 9032 56810
rect 8094 56754 8102 56790
rect 8030 56738 8102 56754
rect 8154 56754 8180 56790
rect 8278 56754 8322 56790
rect 8402 56754 8464 56790
rect 8154 56738 8226 56754
rect 8278 56738 8350 56754
rect 8402 56738 8474 56754
rect 8526 56738 8598 56790
rect 8662 56754 8722 56790
rect 8804 56754 8846 56790
rect 8946 56754 8970 56790
rect 8650 56738 8722 56754
rect 8774 56738 8846 56754
rect 8898 56738 8970 56754
rect 9022 56754 9032 56790
rect 9088 56790 9174 56810
rect 9230 56790 9316 56810
rect 9372 56790 9458 56810
rect 9514 56790 9600 56810
rect 9656 56790 9742 56810
rect 9798 56790 9884 56810
rect 9940 56790 10026 56810
rect 9088 56754 9094 56790
rect 9022 56738 9094 56754
rect 9146 56754 9174 56790
rect 9270 56754 9316 56790
rect 9394 56754 9458 56790
rect 9146 56738 9218 56754
rect 9270 56738 9342 56754
rect 9394 56738 9466 56754
rect 9518 56738 9590 56790
rect 9656 56754 9714 56790
rect 9798 56754 9838 56790
rect 9940 56754 9962 56790
rect 9642 56738 9714 56754
rect 9766 56738 9838 56754
rect 9890 56738 9962 56754
rect 10014 56754 10026 56790
rect 10082 56790 10168 56810
rect 10224 56790 10310 56810
rect 10366 56790 10452 56810
rect 10508 56790 10594 56810
rect 10650 56790 10736 56810
rect 10792 56790 10878 56810
rect 10934 56790 11020 56810
rect 10082 56754 10086 56790
rect 10014 56738 10086 56754
rect 10138 56754 10168 56790
rect 10262 56754 10310 56790
rect 10386 56754 10452 56790
rect 10138 56738 10210 56754
rect 10262 56738 10334 56754
rect 10386 56738 10458 56754
rect 10510 56738 10582 56790
rect 10650 56754 10706 56790
rect 10792 56754 10830 56790
rect 10934 56754 10954 56790
rect 10634 56738 10706 56754
rect 10758 56738 10830 56754
rect 10882 56738 10954 56754
rect 11006 56754 11020 56790
rect 11076 56790 11162 56810
rect 11218 56790 11304 56810
rect 11360 56790 11446 56810
rect 11502 56790 11588 56810
rect 11644 56790 11730 56810
rect 11786 56790 11872 56810
rect 11928 56790 12014 56810
rect 11076 56754 11078 56790
rect 11006 56738 11078 56754
rect 11130 56754 11162 56790
rect 11254 56754 11304 56790
rect 11378 56754 11446 56790
rect 11130 56738 11202 56754
rect 11254 56738 11326 56754
rect 11378 56738 11450 56754
rect 11502 56738 11574 56790
rect 11644 56754 11698 56790
rect 11786 56754 11822 56790
rect 11928 56754 11946 56790
rect 11626 56738 11698 56754
rect 11750 56738 11822 56754
rect 11874 56738 11946 56754
rect 11998 56754 12014 56790
rect 12070 56790 12156 56810
rect 12212 56790 12298 56810
rect 12354 56790 12440 56810
rect 12496 56790 12582 56810
rect 12638 56790 12724 56810
rect 12780 56790 12866 56810
rect 11998 56738 12070 56754
rect 12122 56754 12156 56790
rect 12246 56754 12298 56790
rect 12370 56754 12440 56790
rect 12496 56754 12566 56790
rect 12638 56754 12690 56790
rect 12780 56754 12814 56790
rect 12122 56738 12194 56754
rect 12246 56738 12318 56754
rect 12370 56738 12442 56754
rect 12494 56738 12566 56754
rect 12618 56738 12690 56754
rect 12742 56738 12814 56754
rect 12922 56790 13008 56810
rect 13064 56790 13150 56810
rect 13206 56790 13292 56810
rect 13348 56790 13434 56810
rect 13490 56790 13576 56810
rect 12922 56754 12938 56790
rect 12866 56738 12938 56754
rect 12990 56754 13008 56790
rect 13114 56754 13150 56790
rect 13238 56754 13292 56790
rect 12990 56738 13062 56754
rect 13114 56738 13186 56754
rect 13238 56738 13310 56754
rect 13362 56738 13434 56790
rect 13490 56754 13558 56790
rect 13632 56754 13642 56810
rect 13486 56738 13558 56754
rect 13610 56738 13642 56754
rect 2490 56668 13642 56738
rect 2490 56612 2500 56668
rect 2556 56666 2642 56668
rect 2698 56666 2784 56668
rect 2840 56666 2926 56668
rect 2982 56666 3068 56668
rect 3124 56666 3210 56668
rect 2574 56614 2642 56666
rect 2698 56614 2770 56666
rect 2840 56614 2894 56666
rect 2982 56614 3018 56666
rect 3124 56614 3142 56666
rect 3194 56614 3210 56666
rect 2556 56612 2642 56614
rect 2698 56612 2784 56614
rect 2840 56612 2926 56614
rect 2982 56612 3068 56614
rect 3124 56612 3210 56614
rect 3266 56666 3352 56668
rect 3408 56666 3494 56668
rect 3550 56666 3636 56668
rect 3692 56666 3778 56668
rect 3834 56666 3920 56668
rect 3976 56666 4062 56668
rect 3318 56614 3352 56666
rect 3442 56614 3494 56666
rect 3566 56614 3636 56666
rect 3692 56614 3762 56666
rect 3834 56614 3886 56666
rect 3976 56614 4010 56666
rect 3266 56612 3352 56614
rect 3408 56612 3494 56614
rect 3550 56612 3636 56614
rect 3692 56612 3778 56614
rect 3834 56612 3920 56614
rect 3976 56612 4062 56614
rect 4118 56666 4204 56668
rect 4260 56666 4346 56668
rect 4402 56666 4488 56668
rect 4544 56666 4630 56668
rect 4686 56666 4772 56668
rect 4828 56666 4914 56668
rect 4970 56666 5056 56668
rect 4118 56614 4134 56666
rect 4186 56614 4204 56666
rect 4310 56614 4346 56666
rect 4434 56614 4488 56666
rect 4558 56614 4630 56666
rect 4686 56614 4754 56666
rect 4828 56614 4878 56666
rect 4970 56614 5002 56666
rect 5054 56614 5056 56666
rect 4118 56612 4204 56614
rect 4260 56612 4346 56614
rect 4402 56612 4488 56614
rect 4544 56612 4630 56614
rect 4686 56612 4772 56614
rect 4828 56612 4914 56614
rect 4970 56612 5056 56614
rect 5112 56666 5198 56668
rect 5254 56666 5340 56668
rect 5396 56666 5482 56668
rect 5538 56666 5624 56668
rect 5680 56666 5766 56668
rect 5822 56666 5908 56668
rect 5964 56666 6050 56668
rect 5112 56614 5126 56666
rect 5178 56614 5198 56666
rect 5302 56614 5340 56666
rect 5426 56614 5482 56666
rect 5550 56614 5622 56666
rect 5680 56614 5746 56666
rect 5822 56614 5870 56666
rect 5964 56614 5994 56666
rect 6046 56614 6050 56666
rect 5112 56612 5198 56614
rect 5254 56612 5340 56614
rect 5396 56612 5482 56614
rect 5538 56612 5624 56614
rect 5680 56612 5766 56614
rect 5822 56612 5908 56614
rect 5964 56612 6050 56614
rect 6106 56666 6192 56668
rect 6248 56666 6334 56668
rect 6390 56666 6476 56668
rect 6532 56666 6618 56668
rect 6674 56666 6760 56668
rect 6816 56666 6902 56668
rect 6958 56666 7044 56668
rect 6106 56614 6118 56666
rect 6170 56614 6192 56666
rect 6294 56614 6334 56666
rect 6418 56614 6476 56666
rect 6542 56614 6614 56666
rect 6674 56614 6738 56666
rect 6816 56614 6862 56666
rect 6958 56614 6986 56666
rect 7038 56614 7044 56666
rect 6106 56612 6192 56614
rect 6248 56612 6334 56614
rect 6390 56612 6476 56614
rect 6532 56612 6618 56614
rect 6674 56612 6760 56614
rect 6816 56612 6902 56614
rect 6958 56612 7044 56614
rect 7100 56666 7186 56668
rect 7242 56666 7328 56668
rect 7384 56666 7470 56668
rect 7526 56666 7612 56668
rect 7668 56666 7754 56668
rect 7810 56666 7896 56668
rect 7952 56666 8038 56668
rect 7100 56614 7110 56666
rect 7162 56614 7186 56666
rect 7286 56614 7328 56666
rect 7410 56614 7470 56666
rect 7534 56614 7606 56666
rect 7668 56614 7730 56666
rect 7810 56614 7854 56666
rect 7952 56614 7978 56666
rect 8030 56614 8038 56666
rect 7100 56612 7186 56614
rect 7242 56612 7328 56614
rect 7384 56612 7470 56614
rect 7526 56612 7612 56614
rect 7668 56612 7754 56614
rect 7810 56612 7896 56614
rect 7952 56612 8038 56614
rect 8094 56666 8180 56668
rect 8236 56666 8322 56668
rect 8378 56666 8464 56668
rect 8520 56666 8606 56668
rect 8662 56666 8748 56668
rect 8804 56666 8890 56668
rect 8946 56666 9032 56668
rect 8094 56614 8102 56666
rect 8154 56614 8180 56666
rect 8278 56614 8322 56666
rect 8402 56614 8464 56666
rect 8526 56614 8598 56666
rect 8662 56614 8722 56666
rect 8804 56614 8846 56666
rect 8946 56614 8970 56666
rect 9022 56614 9032 56666
rect 8094 56612 8180 56614
rect 8236 56612 8322 56614
rect 8378 56612 8464 56614
rect 8520 56612 8606 56614
rect 8662 56612 8748 56614
rect 8804 56612 8890 56614
rect 8946 56612 9032 56614
rect 9088 56666 9174 56668
rect 9230 56666 9316 56668
rect 9372 56666 9458 56668
rect 9514 56666 9600 56668
rect 9656 56666 9742 56668
rect 9798 56666 9884 56668
rect 9940 56666 10026 56668
rect 9088 56614 9094 56666
rect 9146 56614 9174 56666
rect 9270 56614 9316 56666
rect 9394 56614 9458 56666
rect 9518 56614 9590 56666
rect 9656 56614 9714 56666
rect 9798 56614 9838 56666
rect 9940 56614 9962 56666
rect 10014 56614 10026 56666
rect 9088 56612 9174 56614
rect 9230 56612 9316 56614
rect 9372 56612 9458 56614
rect 9514 56612 9600 56614
rect 9656 56612 9742 56614
rect 9798 56612 9884 56614
rect 9940 56612 10026 56614
rect 10082 56666 10168 56668
rect 10224 56666 10310 56668
rect 10366 56666 10452 56668
rect 10508 56666 10594 56668
rect 10650 56666 10736 56668
rect 10792 56666 10878 56668
rect 10934 56666 11020 56668
rect 10082 56614 10086 56666
rect 10138 56614 10168 56666
rect 10262 56614 10310 56666
rect 10386 56614 10452 56666
rect 10510 56614 10582 56666
rect 10650 56614 10706 56666
rect 10792 56614 10830 56666
rect 10934 56614 10954 56666
rect 11006 56614 11020 56666
rect 10082 56612 10168 56614
rect 10224 56612 10310 56614
rect 10366 56612 10452 56614
rect 10508 56612 10594 56614
rect 10650 56612 10736 56614
rect 10792 56612 10878 56614
rect 10934 56612 11020 56614
rect 11076 56666 11162 56668
rect 11218 56666 11304 56668
rect 11360 56666 11446 56668
rect 11502 56666 11588 56668
rect 11644 56666 11730 56668
rect 11786 56666 11872 56668
rect 11928 56666 12014 56668
rect 11076 56614 11078 56666
rect 11130 56614 11162 56666
rect 11254 56614 11304 56666
rect 11378 56614 11446 56666
rect 11502 56614 11574 56666
rect 11644 56614 11698 56666
rect 11786 56614 11822 56666
rect 11928 56614 11946 56666
rect 11998 56614 12014 56666
rect 11076 56612 11162 56614
rect 11218 56612 11304 56614
rect 11360 56612 11446 56614
rect 11502 56612 11588 56614
rect 11644 56612 11730 56614
rect 11786 56612 11872 56614
rect 11928 56612 12014 56614
rect 12070 56666 12156 56668
rect 12212 56666 12298 56668
rect 12354 56666 12440 56668
rect 12496 56666 12582 56668
rect 12638 56666 12724 56668
rect 12780 56666 12866 56668
rect 12122 56614 12156 56666
rect 12246 56614 12298 56666
rect 12370 56614 12440 56666
rect 12496 56614 12566 56666
rect 12638 56614 12690 56666
rect 12780 56614 12814 56666
rect 12070 56612 12156 56614
rect 12212 56612 12298 56614
rect 12354 56612 12440 56614
rect 12496 56612 12582 56614
rect 12638 56612 12724 56614
rect 12780 56612 12866 56614
rect 12922 56666 13008 56668
rect 13064 56666 13150 56668
rect 13206 56666 13292 56668
rect 13348 56666 13434 56668
rect 13490 56666 13576 56668
rect 12922 56614 12938 56666
rect 12990 56614 13008 56666
rect 13114 56614 13150 56666
rect 13238 56614 13292 56666
rect 13362 56614 13434 56666
rect 13490 56614 13558 56666
rect 12922 56612 13008 56614
rect 13064 56612 13150 56614
rect 13206 56612 13292 56614
rect 13348 56612 13434 56614
rect 13490 56612 13576 56614
rect 13632 56612 13642 56668
rect 2490 56542 13642 56612
rect 2490 56526 2522 56542
rect 2574 56526 2646 56542
rect 2490 56470 2500 56526
rect 2574 56490 2642 56526
rect 2698 56490 2770 56542
rect 2822 56526 2894 56542
rect 2946 56526 3018 56542
rect 3070 56526 3142 56542
rect 2840 56490 2894 56526
rect 2982 56490 3018 56526
rect 3124 56490 3142 56526
rect 3194 56526 3266 56542
rect 3194 56490 3210 56526
rect 2556 56470 2642 56490
rect 2698 56470 2784 56490
rect 2840 56470 2926 56490
rect 2982 56470 3068 56490
rect 3124 56470 3210 56490
rect 3318 56526 3390 56542
rect 3442 56526 3514 56542
rect 3566 56526 3638 56542
rect 3690 56526 3762 56542
rect 3814 56526 3886 56542
rect 3938 56526 4010 56542
rect 3318 56490 3352 56526
rect 3442 56490 3494 56526
rect 3566 56490 3636 56526
rect 3692 56490 3762 56526
rect 3834 56490 3886 56526
rect 3976 56490 4010 56526
rect 4062 56526 4134 56542
rect 3266 56470 3352 56490
rect 3408 56470 3494 56490
rect 3550 56470 3636 56490
rect 3692 56470 3778 56490
rect 3834 56470 3920 56490
rect 3976 56470 4062 56490
rect 4118 56490 4134 56526
rect 4186 56526 4258 56542
rect 4310 56526 4382 56542
rect 4434 56526 4506 56542
rect 4186 56490 4204 56526
rect 4310 56490 4346 56526
rect 4434 56490 4488 56526
rect 4558 56490 4630 56542
rect 4682 56526 4754 56542
rect 4806 56526 4878 56542
rect 4930 56526 5002 56542
rect 4686 56490 4754 56526
rect 4828 56490 4878 56526
rect 4970 56490 5002 56526
rect 5054 56526 5126 56542
rect 5054 56490 5056 56526
rect 4118 56470 4204 56490
rect 4260 56470 4346 56490
rect 4402 56470 4488 56490
rect 4544 56470 4630 56490
rect 4686 56470 4772 56490
rect 4828 56470 4914 56490
rect 4970 56470 5056 56490
rect 5112 56490 5126 56526
rect 5178 56526 5250 56542
rect 5302 56526 5374 56542
rect 5426 56526 5498 56542
rect 5178 56490 5198 56526
rect 5302 56490 5340 56526
rect 5426 56490 5482 56526
rect 5550 56490 5622 56542
rect 5674 56526 5746 56542
rect 5798 56526 5870 56542
rect 5922 56526 5994 56542
rect 5680 56490 5746 56526
rect 5822 56490 5870 56526
rect 5964 56490 5994 56526
rect 6046 56526 6118 56542
rect 6046 56490 6050 56526
rect 5112 56470 5198 56490
rect 5254 56470 5340 56490
rect 5396 56470 5482 56490
rect 5538 56470 5624 56490
rect 5680 56470 5766 56490
rect 5822 56470 5908 56490
rect 5964 56470 6050 56490
rect 6106 56490 6118 56526
rect 6170 56526 6242 56542
rect 6294 56526 6366 56542
rect 6418 56526 6490 56542
rect 6170 56490 6192 56526
rect 6294 56490 6334 56526
rect 6418 56490 6476 56526
rect 6542 56490 6614 56542
rect 6666 56526 6738 56542
rect 6790 56526 6862 56542
rect 6914 56526 6986 56542
rect 6674 56490 6738 56526
rect 6816 56490 6862 56526
rect 6958 56490 6986 56526
rect 7038 56526 7110 56542
rect 7038 56490 7044 56526
rect 6106 56470 6192 56490
rect 6248 56470 6334 56490
rect 6390 56470 6476 56490
rect 6532 56470 6618 56490
rect 6674 56470 6760 56490
rect 6816 56470 6902 56490
rect 6958 56470 7044 56490
rect 7100 56490 7110 56526
rect 7162 56526 7234 56542
rect 7286 56526 7358 56542
rect 7410 56526 7482 56542
rect 7162 56490 7186 56526
rect 7286 56490 7328 56526
rect 7410 56490 7470 56526
rect 7534 56490 7606 56542
rect 7658 56526 7730 56542
rect 7782 56526 7854 56542
rect 7906 56526 7978 56542
rect 7668 56490 7730 56526
rect 7810 56490 7854 56526
rect 7952 56490 7978 56526
rect 8030 56526 8102 56542
rect 8030 56490 8038 56526
rect 7100 56470 7186 56490
rect 7242 56470 7328 56490
rect 7384 56470 7470 56490
rect 7526 56470 7612 56490
rect 7668 56470 7754 56490
rect 7810 56470 7896 56490
rect 7952 56470 8038 56490
rect 8094 56490 8102 56526
rect 8154 56526 8226 56542
rect 8278 56526 8350 56542
rect 8402 56526 8474 56542
rect 8154 56490 8180 56526
rect 8278 56490 8322 56526
rect 8402 56490 8464 56526
rect 8526 56490 8598 56542
rect 8650 56526 8722 56542
rect 8774 56526 8846 56542
rect 8898 56526 8970 56542
rect 8662 56490 8722 56526
rect 8804 56490 8846 56526
rect 8946 56490 8970 56526
rect 9022 56526 9094 56542
rect 9022 56490 9032 56526
rect 8094 56470 8180 56490
rect 8236 56470 8322 56490
rect 8378 56470 8464 56490
rect 8520 56470 8606 56490
rect 8662 56470 8748 56490
rect 8804 56470 8890 56490
rect 8946 56470 9032 56490
rect 9088 56490 9094 56526
rect 9146 56526 9218 56542
rect 9270 56526 9342 56542
rect 9394 56526 9466 56542
rect 9146 56490 9174 56526
rect 9270 56490 9316 56526
rect 9394 56490 9458 56526
rect 9518 56490 9590 56542
rect 9642 56526 9714 56542
rect 9766 56526 9838 56542
rect 9890 56526 9962 56542
rect 9656 56490 9714 56526
rect 9798 56490 9838 56526
rect 9940 56490 9962 56526
rect 10014 56526 10086 56542
rect 10014 56490 10026 56526
rect 9088 56470 9174 56490
rect 9230 56470 9316 56490
rect 9372 56470 9458 56490
rect 9514 56470 9600 56490
rect 9656 56470 9742 56490
rect 9798 56470 9884 56490
rect 9940 56470 10026 56490
rect 10082 56490 10086 56526
rect 10138 56526 10210 56542
rect 10262 56526 10334 56542
rect 10386 56526 10458 56542
rect 10138 56490 10168 56526
rect 10262 56490 10310 56526
rect 10386 56490 10452 56526
rect 10510 56490 10582 56542
rect 10634 56526 10706 56542
rect 10758 56526 10830 56542
rect 10882 56526 10954 56542
rect 10650 56490 10706 56526
rect 10792 56490 10830 56526
rect 10934 56490 10954 56526
rect 11006 56526 11078 56542
rect 11006 56490 11020 56526
rect 10082 56470 10168 56490
rect 10224 56470 10310 56490
rect 10366 56470 10452 56490
rect 10508 56470 10594 56490
rect 10650 56470 10736 56490
rect 10792 56470 10878 56490
rect 10934 56470 11020 56490
rect 11076 56490 11078 56526
rect 11130 56526 11202 56542
rect 11254 56526 11326 56542
rect 11378 56526 11450 56542
rect 11130 56490 11162 56526
rect 11254 56490 11304 56526
rect 11378 56490 11446 56526
rect 11502 56490 11574 56542
rect 11626 56526 11698 56542
rect 11750 56526 11822 56542
rect 11874 56526 11946 56542
rect 11644 56490 11698 56526
rect 11786 56490 11822 56526
rect 11928 56490 11946 56526
rect 11998 56526 12070 56542
rect 11998 56490 12014 56526
rect 11076 56470 11162 56490
rect 11218 56470 11304 56490
rect 11360 56470 11446 56490
rect 11502 56470 11588 56490
rect 11644 56470 11730 56490
rect 11786 56470 11872 56490
rect 11928 56470 12014 56490
rect 12122 56526 12194 56542
rect 12246 56526 12318 56542
rect 12370 56526 12442 56542
rect 12494 56526 12566 56542
rect 12618 56526 12690 56542
rect 12742 56526 12814 56542
rect 12122 56490 12156 56526
rect 12246 56490 12298 56526
rect 12370 56490 12440 56526
rect 12496 56490 12566 56526
rect 12638 56490 12690 56526
rect 12780 56490 12814 56526
rect 12866 56526 12938 56542
rect 12070 56470 12156 56490
rect 12212 56470 12298 56490
rect 12354 56470 12440 56490
rect 12496 56470 12582 56490
rect 12638 56470 12724 56490
rect 12780 56470 12866 56490
rect 12922 56490 12938 56526
rect 12990 56526 13062 56542
rect 13114 56526 13186 56542
rect 13238 56526 13310 56542
rect 12990 56490 13008 56526
rect 13114 56490 13150 56526
rect 13238 56490 13292 56526
rect 13362 56490 13434 56542
rect 13486 56526 13558 56542
rect 13610 56526 13642 56542
rect 13490 56490 13558 56526
rect 12922 56470 13008 56490
rect 13064 56470 13150 56490
rect 13206 56470 13292 56490
rect 13348 56470 13434 56490
rect 13490 56470 13576 56490
rect 13632 56470 13642 56526
rect 2490 56460 13642 56470
rect 2670 56345 13350 56377
rect 2670 56189 2682 56345
rect 2838 56189 3682 56345
rect 3838 56189 4182 56345
rect 4338 56189 5182 56345
rect 5338 56189 5682 56345
rect 5838 56189 6682 56345
rect 6838 56189 7182 56345
rect 7338 56189 8182 56345
rect 8338 56189 8682 56345
rect 8838 56189 9682 56345
rect 9838 56189 10182 56345
rect 10338 56189 11182 56345
rect 11338 56189 11682 56345
rect 11838 56189 12682 56345
rect 12838 56189 13182 56345
rect 13338 56189 13350 56345
rect 2670 56161 13350 56189
rect 2490 56068 13642 56078
rect 2490 56012 2500 56068
rect 2556 56048 2642 56068
rect 2698 56048 2784 56068
rect 2840 56048 2926 56068
rect 2982 56048 3068 56068
rect 3124 56048 3210 56068
rect 2574 56012 2642 56048
rect 2490 55996 2522 56012
rect 2574 55996 2646 56012
rect 2698 55996 2770 56048
rect 2840 56012 2894 56048
rect 2982 56012 3018 56048
rect 3124 56012 3142 56048
rect 2822 55996 2894 56012
rect 2946 55996 3018 56012
rect 3070 55996 3142 56012
rect 3194 56012 3210 56048
rect 3266 56048 3352 56068
rect 3408 56048 3494 56068
rect 3550 56048 3636 56068
rect 3692 56048 3778 56068
rect 3834 56048 3920 56068
rect 3976 56048 4062 56068
rect 3194 55996 3266 56012
rect 3318 56012 3352 56048
rect 3442 56012 3494 56048
rect 3566 56012 3636 56048
rect 3692 56012 3762 56048
rect 3834 56012 3886 56048
rect 3976 56012 4010 56048
rect 3318 55996 3390 56012
rect 3442 55996 3514 56012
rect 3566 55996 3638 56012
rect 3690 55996 3762 56012
rect 3814 55996 3886 56012
rect 3938 55996 4010 56012
rect 4118 56048 4204 56068
rect 4260 56048 4346 56068
rect 4402 56048 4488 56068
rect 4544 56048 4630 56068
rect 4686 56048 4772 56068
rect 4828 56048 4914 56068
rect 4970 56048 5056 56068
rect 4118 56012 4134 56048
rect 4062 55996 4134 56012
rect 4186 56012 4204 56048
rect 4310 56012 4346 56048
rect 4434 56012 4488 56048
rect 4186 55996 4258 56012
rect 4310 55996 4382 56012
rect 4434 55996 4506 56012
rect 4558 55996 4630 56048
rect 4686 56012 4754 56048
rect 4828 56012 4878 56048
rect 4970 56012 5002 56048
rect 4682 55996 4754 56012
rect 4806 55996 4878 56012
rect 4930 55996 5002 56012
rect 5054 56012 5056 56048
rect 5112 56048 5198 56068
rect 5254 56048 5340 56068
rect 5396 56048 5482 56068
rect 5538 56048 5624 56068
rect 5680 56048 5766 56068
rect 5822 56048 5908 56068
rect 5964 56048 6050 56068
rect 5112 56012 5126 56048
rect 5054 55996 5126 56012
rect 5178 56012 5198 56048
rect 5302 56012 5340 56048
rect 5426 56012 5482 56048
rect 5178 55996 5250 56012
rect 5302 55996 5374 56012
rect 5426 55996 5498 56012
rect 5550 55996 5622 56048
rect 5680 56012 5746 56048
rect 5822 56012 5870 56048
rect 5964 56012 5994 56048
rect 5674 55996 5746 56012
rect 5798 55996 5870 56012
rect 5922 55996 5994 56012
rect 6046 56012 6050 56048
rect 6106 56048 6192 56068
rect 6248 56048 6334 56068
rect 6390 56048 6476 56068
rect 6532 56048 6618 56068
rect 6674 56048 6760 56068
rect 6816 56048 6902 56068
rect 6958 56048 7044 56068
rect 6106 56012 6118 56048
rect 6046 55996 6118 56012
rect 6170 56012 6192 56048
rect 6294 56012 6334 56048
rect 6418 56012 6476 56048
rect 6170 55996 6242 56012
rect 6294 55996 6366 56012
rect 6418 55996 6490 56012
rect 6542 55996 6614 56048
rect 6674 56012 6738 56048
rect 6816 56012 6862 56048
rect 6958 56012 6986 56048
rect 6666 55996 6738 56012
rect 6790 55996 6862 56012
rect 6914 55996 6986 56012
rect 7038 56012 7044 56048
rect 7100 56048 7186 56068
rect 7242 56048 7328 56068
rect 7384 56048 7470 56068
rect 7526 56048 7612 56068
rect 7668 56048 7754 56068
rect 7810 56048 7896 56068
rect 7952 56048 8038 56068
rect 7100 56012 7110 56048
rect 7038 55996 7110 56012
rect 7162 56012 7186 56048
rect 7286 56012 7328 56048
rect 7410 56012 7470 56048
rect 7162 55996 7234 56012
rect 7286 55996 7358 56012
rect 7410 55996 7482 56012
rect 7534 55996 7606 56048
rect 7668 56012 7730 56048
rect 7810 56012 7854 56048
rect 7952 56012 7978 56048
rect 7658 55996 7730 56012
rect 7782 55996 7854 56012
rect 7906 55996 7978 56012
rect 8030 56012 8038 56048
rect 8094 56048 8180 56068
rect 8236 56048 8322 56068
rect 8378 56048 8464 56068
rect 8520 56048 8606 56068
rect 8662 56048 8748 56068
rect 8804 56048 8890 56068
rect 8946 56048 9032 56068
rect 8094 56012 8102 56048
rect 8030 55996 8102 56012
rect 8154 56012 8180 56048
rect 8278 56012 8322 56048
rect 8402 56012 8464 56048
rect 8154 55996 8226 56012
rect 8278 55996 8350 56012
rect 8402 55996 8474 56012
rect 8526 55996 8598 56048
rect 8662 56012 8722 56048
rect 8804 56012 8846 56048
rect 8946 56012 8970 56048
rect 8650 55996 8722 56012
rect 8774 55996 8846 56012
rect 8898 55996 8970 56012
rect 9022 56012 9032 56048
rect 9088 56048 9174 56068
rect 9230 56048 9316 56068
rect 9372 56048 9458 56068
rect 9514 56048 9600 56068
rect 9656 56048 9742 56068
rect 9798 56048 9884 56068
rect 9940 56048 10026 56068
rect 9088 56012 9094 56048
rect 9022 55996 9094 56012
rect 9146 56012 9174 56048
rect 9270 56012 9316 56048
rect 9394 56012 9458 56048
rect 9146 55996 9218 56012
rect 9270 55996 9342 56012
rect 9394 55996 9466 56012
rect 9518 55996 9590 56048
rect 9656 56012 9714 56048
rect 9798 56012 9838 56048
rect 9940 56012 9962 56048
rect 9642 55996 9714 56012
rect 9766 55996 9838 56012
rect 9890 55996 9962 56012
rect 10014 56012 10026 56048
rect 10082 56048 10168 56068
rect 10224 56048 10310 56068
rect 10366 56048 10452 56068
rect 10508 56048 10594 56068
rect 10650 56048 10736 56068
rect 10792 56048 10878 56068
rect 10934 56048 11020 56068
rect 10082 56012 10086 56048
rect 10014 55996 10086 56012
rect 10138 56012 10168 56048
rect 10262 56012 10310 56048
rect 10386 56012 10452 56048
rect 10138 55996 10210 56012
rect 10262 55996 10334 56012
rect 10386 55996 10458 56012
rect 10510 55996 10582 56048
rect 10650 56012 10706 56048
rect 10792 56012 10830 56048
rect 10934 56012 10954 56048
rect 10634 55996 10706 56012
rect 10758 55996 10830 56012
rect 10882 55996 10954 56012
rect 11006 56012 11020 56048
rect 11076 56048 11162 56068
rect 11218 56048 11304 56068
rect 11360 56048 11446 56068
rect 11502 56048 11588 56068
rect 11644 56048 11730 56068
rect 11786 56048 11872 56068
rect 11928 56048 12014 56068
rect 11076 56012 11078 56048
rect 11006 55996 11078 56012
rect 11130 56012 11162 56048
rect 11254 56012 11304 56048
rect 11378 56012 11446 56048
rect 11130 55996 11202 56012
rect 11254 55996 11326 56012
rect 11378 55996 11450 56012
rect 11502 55996 11574 56048
rect 11644 56012 11698 56048
rect 11786 56012 11822 56048
rect 11928 56012 11946 56048
rect 11626 55996 11698 56012
rect 11750 55996 11822 56012
rect 11874 55996 11946 56012
rect 11998 56012 12014 56048
rect 12070 56048 12156 56068
rect 12212 56048 12298 56068
rect 12354 56048 12440 56068
rect 12496 56048 12582 56068
rect 12638 56048 12724 56068
rect 12780 56048 12866 56068
rect 11998 55996 12070 56012
rect 12122 56012 12156 56048
rect 12246 56012 12298 56048
rect 12370 56012 12440 56048
rect 12496 56012 12566 56048
rect 12638 56012 12690 56048
rect 12780 56012 12814 56048
rect 12122 55996 12194 56012
rect 12246 55996 12318 56012
rect 12370 55996 12442 56012
rect 12494 55996 12566 56012
rect 12618 55996 12690 56012
rect 12742 55996 12814 56012
rect 12922 56048 13008 56068
rect 13064 56048 13150 56068
rect 13206 56048 13292 56068
rect 13348 56048 13434 56068
rect 13490 56048 13576 56068
rect 12922 56012 12938 56048
rect 12866 55996 12938 56012
rect 12990 56012 13008 56048
rect 13114 56012 13150 56048
rect 13238 56012 13292 56048
rect 12990 55996 13062 56012
rect 13114 55996 13186 56012
rect 13238 55996 13310 56012
rect 13362 55996 13434 56048
rect 13490 56012 13558 56048
rect 13632 56012 13642 56068
rect 13486 55996 13558 56012
rect 13610 55996 13642 56012
rect 2490 55926 13642 55996
rect 2490 55870 2500 55926
rect 2556 55924 2642 55926
rect 2698 55924 2784 55926
rect 2840 55924 2926 55926
rect 2982 55924 3068 55926
rect 3124 55924 3210 55926
rect 2574 55872 2642 55924
rect 2698 55872 2770 55924
rect 2840 55872 2894 55924
rect 2982 55872 3018 55924
rect 3124 55872 3142 55924
rect 3194 55872 3210 55924
rect 2556 55870 2642 55872
rect 2698 55870 2784 55872
rect 2840 55870 2926 55872
rect 2982 55870 3068 55872
rect 3124 55870 3210 55872
rect 3266 55924 3352 55926
rect 3408 55924 3494 55926
rect 3550 55924 3636 55926
rect 3692 55924 3778 55926
rect 3834 55924 3920 55926
rect 3976 55924 4062 55926
rect 3318 55872 3352 55924
rect 3442 55872 3494 55924
rect 3566 55872 3636 55924
rect 3692 55872 3762 55924
rect 3834 55872 3886 55924
rect 3976 55872 4010 55924
rect 3266 55870 3352 55872
rect 3408 55870 3494 55872
rect 3550 55870 3636 55872
rect 3692 55870 3778 55872
rect 3834 55870 3920 55872
rect 3976 55870 4062 55872
rect 4118 55924 4204 55926
rect 4260 55924 4346 55926
rect 4402 55924 4488 55926
rect 4544 55924 4630 55926
rect 4686 55924 4772 55926
rect 4828 55924 4914 55926
rect 4970 55924 5056 55926
rect 4118 55872 4134 55924
rect 4186 55872 4204 55924
rect 4310 55872 4346 55924
rect 4434 55872 4488 55924
rect 4558 55872 4630 55924
rect 4686 55872 4754 55924
rect 4828 55872 4878 55924
rect 4970 55872 5002 55924
rect 5054 55872 5056 55924
rect 4118 55870 4204 55872
rect 4260 55870 4346 55872
rect 4402 55870 4488 55872
rect 4544 55870 4630 55872
rect 4686 55870 4772 55872
rect 4828 55870 4914 55872
rect 4970 55870 5056 55872
rect 5112 55924 5198 55926
rect 5254 55924 5340 55926
rect 5396 55924 5482 55926
rect 5538 55924 5624 55926
rect 5680 55924 5766 55926
rect 5822 55924 5908 55926
rect 5964 55924 6050 55926
rect 5112 55872 5126 55924
rect 5178 55872 5198 55924
rect 5302 55872 5340 55924
rect 5426 55872 5482 55924
rect 5550 55872 5622 55924
rect 5680 55872 5746 55924
rect 5822 55872 5870 55924
rect 5964 55872 5994 55924
rect 6046 55872 6050 55924
rect 5112 55870 5198 55872
rect 5254 55870 5340 55872
rect 5396 55870 5482 55872
rect 5538 55870 5624 55872
rect 5680 55870 5766 55872
rect 5822 55870 5908 55872
rect 5964 55870 6050 55872
rect 6106 55924 6192 55926
rect 6248 55924 6334 55926
rect 6390 55924 6476 55926
rect 6532 55924 6618 55926
rect 6674 55924 6760 55926
rect 6816 55924 6902 55926
rect 6958 55924 7044 55926
rect 6106 55872 6118 55924
rect 6170 55872 6192 55924
rect 6294 55872 6334 55924
rect 6418 55872 6476 55924
rect 6542 55872 6614 55924
rect 6674 55872 6738 55924
rect 6816 55872 6862 55924
rect 6958 55872 6986 55924
rect 7038 55872 7044 55924
rect 6106 55870 6192 55872
rect 6248 55870 6334 55872
rect 6390 55870 6476 55872
rect 6532 55870 6618 55872
rect 6674 55870 6760 55872
rect 6816 55870 6902 55872
rect 6958 55870 7044 55872
rect 7100 55924 7186 55926
rect 7242 55924 7328 55926
rect 7384 55924 7470 55926
rect 7526 55924 7612 55926
rect 7668 55924 7754 55926
rect 7810 55924 7896 55926
rect 7952 55924 8038 55926
rect 7100 55872 7110 55924
rect 7162 55872 7186 55924
rect 7286 55872 7328 55924
rect 7410 55872 7470 55924
rect 7534 55872 7606 55924
rect 7668 55872 7730 55924
rect 7810 55872 7854 55924
rect 7952 55872 7978 55924
rect 8030 55872 8038 55924
rect 7100 55870 7186 55872
rect 7242 55870 7328 55872
rect 7384 55870 7470 55872
rect 7526 55870 7612 55872
rect 7668 55870 7754 55872
rect 7810 55870 7896 55872
rect 7952 55870 8038 55872
rect 8094 55924 8180 55926
rect 8236 55924 8322 55926
rect 8378 55924 8464 55926
rect 8520 55924 8606 55926
rect 8662 55924 8748 55926
rect 8804 55924 8890 55926
rect 8946 55924 9032 55926
rect 8094 55872 8102 55924
rect 8154 55872 8180 55924
rect 8278 55872 8322 55924
rect 8402 55872 8464 55924
rect 8526 55872 8598 55924
rect 8662 55872 8722 55924
rect 8804 55872 8846 55924
rect 8946 55872 8970 55924
rect 9022 55872 9032 55924
rect 8094 55870 8180 55872
rect 8236 55870 8322 55872
rect 8378 55870 8464 55872
rect 8520 55870 8606 55872
rect 8662 55870 8748 55872
rect 8804 55870 8890 55872
rect 8946 55870 9032 55872
rect 9088 55924 9174 55926
rect 9230 55924 9316 55926
rect 9372 55924 9458 55926
rect 9514 55924 9600 55926
rect 9656 55924 9742 55926
rect 9798 55924 9884 55926
rect 9940 55924 10026 55926
rect 9088 55872 9094 55924
rect 9146 55872 9174 55924
rect 9270 55872 9316 55924
rect 9394 55872 9458 55924
rect 9518 55872 9590 55924
rect 9656 55872 9714 55924
rect 9798 55872 9838 55924
rect 9940 55872 9962 55924
rect 10014 55872 10026 55924
rect 9088 55870 9174 55872
rect 9230 55870 9316 55872
rect 9372 55870 9458 55872
rect 9514 55870 9600 55872
rect 9656 55870 9742 55872
rect 9798 55870 9884 55872
rect 9940 55870 10026 55872
rect 10082 55924 10168 55926
rect 10224 55924 10310 55926
rect 10366 55924 10452 55926
rect 10508 55924 10594 55926
rect 10650 55924 10736 55926
rect 10792 55924 10878 55926
rect 10934 55924 11020 55926
rect 10082 55872 10086 55924
rect 10138 55872 10168 55924
rect 10262 55872 10310 55924
rect 10386 55872 10452 55924
rect 10510 55872 10582 55924
rect 10650 55872 10706 55924
rect 10792 55872 10830 55924
rect 10934 55872 10954 55924
rect 11006 55872 11020 55924
rect 10082 55870 10168 55872
rect 10224 55870 10310 55872
rect 10366 55870 10452 55872
rect 10508 55870 10594 55872
rect 10650 55870 10736 55872
rect 10792 55870 10878 55872
rect 10934 55870 11020 55872
rect 11076 55924 11162 55926
rect 11218 55924 11304 55926
rect 11360 55924 11446 55926
rect 11502 55924 11588 55926
rect 11644 55924 11730 55926
rect 11786 55924 11872 55926
rect 11928 55924 12014 55926
rect 11076 55872 11078 55924
rect 11130 55872 11162 55924
rect 11254 55872 11304 55924
rect 11378 55872 11446 55924
rect 11502 55872 11574 55924
rect 11644 55872 11698 55924
rect 11786 55872 11822 55924
rect 11928 55872 11946 55924
rect 11998 55872 12014 55924
rect 11076 55870 11162 55872
rect 11218 55870 11304 55872
rect 11360 55870 11446 55872
rect 11502 55870 11588 55872
rect 11644 55870 11730 55872
rect 11786 55870 11872 55872
rect 11928 55870 12014 55872
rect 12070 55924 12156 55926
rect 12212 55924 12298 55926
rect 12354 55924 12440 55926
rect 12496 55924 12582 55926
rect 12638 55924 12724 55926
rect 12780 55924 12866 55926
rect 12122 55872 12156 55924
rect 12246 55872 12298 55924
rect 12370 55872 12440 55924
rect 12496 55872 12566 55924
rect 12638 55872 12690 55924
rect 12780 55872 12814 55924
rect 12070 55870 12156 55872
rect 12212 55870 12298 55872
rect 12354 55870 12440 55872
rect 12496 55870 12582 55872
rect 12638 55870 12724 55872
rect 12780 55870 12866 55872
rect 12922 55924 13008 55926
rect 13064 55924 13150 55926
rect 13206 55924 13292 55926
rect 13348 55924 13434 55926
rect 13490 55924 13576 55926
rect 12922 55872 12938 55924
rect 12990 55872 13008 55924
rect 13114 55872 13150 55924
rect 13238 55872 13292 55924
rect 13362 55872 13434 55924
rect 13490 55872 13558 55924
rect 12922 55870 13008 55872
rect 13064 55870 13150 55872
rect 13206 55870 13292 55872
rect 13348 55870 13434 55872
rect 13490 55870 13576 55872
rect 13632 55870 13642 55926
rect 2490 55800 13642 55870
rect 2490 55784 2522 55800
rect 2574 55784 2646 55800
rect 2490 55728 2500 55784
rect 2574 55748 2642 55784
rect 2698 55748 2770 55800
rect 2822 55784 2894 55800
rect 2946 55784 3018 55800
rect 3070 55784 3142 55800
rect 2840 55748 2894 55784
rect 2982 55748 3018 55784
rect 3124 55748 3142 55784
rect 3194 55784 3266 55800
rect 3194 55748 3210 55784
rect 2556 55728 2642 55748
rect 2698 55728 2784 55748
rect 2840 55728 2926 55748
rect 2982 55728 3068 55748
rect 3124 55728 3210 55748
rect 3318 55784 3390 55800
rect 3442 55784 3514 55800
rect 3566 55784 3638 55800
rect 3690 55784 3762 55800
rect 3814 55784 3886 55800
rect 3938 55784 4010 55800
rect 3318 55748 3352 55784
rect 3442 55748 3494 55784
rect 3566 55748 3636 55784
rect 3692 55748 3762 55784
rect 3834 55748 3886 55784
rect 3976 55748 4010 55784
rect 4062 55784 4134 55800
rect 3266 55728 3352 55748
rect 3408 55728 3494 55748
rect 3550 55728 3636 55748
rect 3692 55728 3778 55748
rect 3834 55728 3920 55748
rect 3976 55728 4062 55748
rect 4118 55748 4134 55784
rect 4186 55784 4258 55800
rect 4310 55784 4382 55800
rect 4434 55784 4506 55800
rect 4186 55748 4204 55784
rect 4310 55748 4346 55784
rect 4434 55748 4488 55784
rect 4558 55748 4630 55800
rect 4682 55784 4754 55800
rect 4806 55784 4878 55800
rect 4930 55784 5002 55800
rect 4686 55748 4754 55784
rect 4828 55748 4878 55784
rect 4970 55748 5002 55784
rect 5054 55784 5126 55800
rect 5054 55748 5056 55784
rect 4118 55728 4204 55748
rect 4260 55728 4346 55748
rect 4402 55728 4488 55748
rect 4544 55728 4630 55748
rect 4686 55728 4772 55748
rect 4828 55728 4914 55748
rect 4970 55728 5056 55748
rect 5112 55748 5126 55784
rect 5178 55784 5250 55800
rect 5302 55784 5374 55800
rect 5426 55784 5498 55800
rect 5178 55748 5198 55784
rect 5302 55748 5340 55784
rect 5426 55748 5482 55784
rect 5550 55748 5622 55800
rect 5674 55784 5746 55800
rect 5798 55784 5870 55800
rect 5922 55784 5994 55800
rect 5680 55748 5746 55784
rect 5822 55748 5870 55784
rect 5964 55748 5994 55784
rect 6046 55784 6118 55800
rect 6046 55748 6050 55784
rect 5112 55728 5198 55748
rect 5254 55728 5340 55748
rect 5396 55728 5482 55748
rect 5538 55728 5624 55748
rect 5680 55728 5766 55748
rect 5822 55728 5908 55748
rect 5964 55728 6050 55748
rect 6106 55748 6118 55784
rect 6170 55784 6242 55800
rect 6294 55784 6366 55800
rect 6418 55784 6490 55800
rect 6170 55748 6192 55784
rect 6294 55748 6334 55784
rect 6418 55748 6476 55784
rect 6542 55748 6614 55800
rect 6666 55784 6738 55800
rect 6790 55784 6862 55800
rect 6914 55784 6986 55800
rect 6674 55748 6738 55784
rect 6816 55748 6862 55784
rect 6958 55748 6986 55784
rect 7038 55784 7110 55800
rect 7038 55748 7044 55784
rect 6106 55728 6192 55748
rect 6248 55728 6334 55748
rect 6390 55728 6476 55748
rect 6532 55728 6618 55748
rect 6674 55728 6760 55748
rect 6816 55728 6902 55748
rect 6958 55728 7044 55748
rect 7100 55748 7110 55784
rect 7162 55784 7234 55800
rect 7286 55784 7358 55800
rect 7410 55784 7482 55800
rect 7162 55748 7186 55784
rect 7286 55748 7328 55784
rect 7410 55748 7470 55784
rect 7534 55748 7606 55800
rect 7658 55784 7730 55800
rect 7782 55784 7854 55800
rect 7906 55784 7978 55800
rect 7668 55748 7730 55784
rect 7810 55748 7854 55784
rect 7952 55748 7978 55784
rect 8030 55784 8102 55800
rect 8030 55748 8038 55784
rect 7100 55728 7186 55748
rect 7242 55728 7328 55748
rect 7384 55728 7470 55748
rect 7526 55728 7612 55748
rect 7668 55728 7754 55748
rect 7810 55728 7896 55748
rect 7952 55728 8038 55748
rect 8094 55748 8102 55784
rect 8154 55784 8226 55800
rect 8278 55784 8350 55800
rect 8402 55784 8474 55800
rect 8154 55748 8180 55784
rect 8278 55748 8322 55784
rect 8402 55748 8464 55784
rect 8526 55748 8598 55800
rect 8650 55784 8722 55800
rect 8774 55784 8846 55800
rect 8898 55784 8970 55800
rect 8662 55748 8722 55784
rect 8804 55748 8846 55784
rect 8946 55748 8970 55784
rect 9022 55784 9094 55800
rect 9022 55748 9032 55784
rect 8094 55728 8180 55748
rect 8236 55728 8322 55748
rect 8378 55728 8464 55748
rect 8520 55728 8606 55748
rect 8662 55728 8748 55748
rect 8804 55728 8890 55748
rect 8946 55728 9032 55748
rect 9088 55748 9094 55784
rect 9146 55784 9218 55800
rect 9270 55784 9342 55800
rect 9394 55784 9466 55800
rect 9146 55748 9174 55784
rect 9270 55748 9316 55784
rect 9394 55748 9458 55784
rect 9518 55748 9590 55800
rect 9642 55784 9714 55800
rect 9766 55784 9838 55800
rect 9890 55784 9962 55800
rect 9656 55748 9714 55784
rect 9798 55748 9838 55784
rect 9940 55748 9962 55784
rect 10014 55784 10086 55800
rect 10014 55748 10026 55784
rect 9088 55728 9174 55748
rect 9230 55728 9316 55748
rect 9372 55728 9458 55748
rect 9514 55728 9600 55748
rect 9656 55728 9742 55748
rect 9798 55728 9884 55748
rect 9940 55728 10026 55748
rect 10082 55748 10086 55784
rect 10138 55784 10210 55800
rect 10262 55784 10334 55800
rect 10386 55784 10458 55800
rect 10138 55748 10168 55784
rect 10262 55748 10310 55784
rect 10386 55748 10452 55784
rect 10510 55748 10582 55800
rect 10634 55784 10706 55800
rect 10758 55784 10830 55800
rect 10882 55784 10954 55800
rect 10650 55748 10706 55784
rect 10792 55748 10830 55784
rect 10934 55748 10954 55784
rect 11006 55784 11078 55800
rect 11006 55748 11020 55784
rect 10082 55728 10168 55748
rect 10224 55728 10310 55748
rect 10366 55728 10452 55748
rect 10508 55728 10594 55748
rect 10650 55728 10736 55748
rect 10792 55728 10878 55748
rect 10934 55728 11020 55748
rect 11076 55748 11078 55784
rect 11130 55784 11202 55800
rect 11254 55784 11326 55800
rect 11378 55784 11450 55800
rect 11130 55748 11162 55784
rect 11254 55748 11304 55784
rect 11378 55748 11446 55784
rect 11502 55748 11574 55800
rect 11626 55784 11698 55800
rect 11750 55784 11822 55800
rect 11874 55784 11946 55800
rect 11644 55748 11698 55784
rect 11786 55748 11822 55784
rect 11928 55748 11946 55784
rect 11998 55784 12070 55800
rect 11998 55748 12014 55784
rect 11076 55728 11162 55748
rect 11218 55728 11304 55748
rect 11360 55728 11446 55748
rect 11502 55728 11588 55748
rect 11644 55728 11730 55748
rect 11786 55728 11872 55748
rect 11928 55728 12014 55748
rect 12122 55784 12194 55800
rect 12246 55784 12318 55800
rect 12370 55784 12442 55800
rect 12494 55784 12566 55800
rect 12618 55784 12690 55800
rect 12742 55784 12814 55800
rect 12122 55748 12156 55784
rect 12246 55748 12298 55784
rect 12370 55748 12440 55784
rect 12496 55748 12566 55784
rect 12638 55748 12690 55784
rect 12780 55748 12814 55784
rect 12866 55784 12938 55800
rect 12070 55728 12156 55748
rect 12212 55728 12298 55748
rect 12354 55728 12440 55748
rect 12496 55728 12582 55748
rect 12638 55728 12724 55748
rect 12780 55728 12866 55748
rect 12922 55748 12938 55784
rect 12990 55784 13062 55800
rect 13114 55784 13186 55800
rect 13238 55784 13310 55800
rect 12990 55748 13008 55784
rect 13114 55748 13150 55784
rect 13238 55748 13292 55784
rect 13362 55748 13434 55800
rect 13486 55784 13558 55800
rect 13610 55784 13642 55800
rect 13490 55748 13558 55784
rect 12922 55728 13008 55748
rect 13064 55728 13150 55748
rect 13206 55728 13292 55748
rect 13348 55728 13434 55748
rect 13490 55728 13576 55748
rect 13632 55728 13642 55784
rect 2490 55718 13642 55728
rect 3470 55479 13350 55555
rect 3470 55459 3546 55479
rect 3470 54471 3482 55459
rect 3534 54471 3546 55459
rect 3470 54459 3546 54471
rect 3693 55459 3769 55479
rect 3693 54471 3705 55459
rect 3757 54471 3769 55459
rect 3693 54459 3769 54471
rect 4162 55459 4238 55479
rect 4162 54471 4174 55459
rect 4226 54471 4238 55459
rect 8030 55459 8106 55479
rect 4758 55404 4834 55416
rect 4758 55397 4770 55404
rect 4822 55397 4834 55404
rect 4758 55341 4768 55397
rect 4824 55341 4834 55397
rect 4758 55255 4770 55341
rect 4822 55255 4834 55341
rect 4758 55199 4768 55255
rect 4824 55199 4834 55255
rect 4758 55113 4770 55199
rect 4822 55113 4834 55199
rect 4758 55057 4768 55113
rect 4824 55057 4834 55113
rect 4758 54971 4770 55057
rect 4822 54971 4834 55057
rect 4758 54915 4768 54971
rect 4824 54915 4834 54971
rect 4758 54829 4770 54915
rect 4822 54829 4834 54915
rect 4758 54773 4768 54829
rect 4824 54773 4834 54829
rect 4758 54687 4770 54773
rect 4822 54687 4834 54773
rect 4758 54631 4768 54687
rect 4824 54631 4834 54687
rect 4758 54624 4770 54631
rect 4822 54624 4834 54631
rect 4758 54612 4834 54624
rect 4938 55404 5014 55416
rect 4938 55397 4950 55404
rect 5002 55397 5014 55404
rect 4938 55341 4948 55397
rect 5004 55341 5014 55397
rect 4938 55255 4950 55341
rect 5002 55255 5014 55341
rect 4938 55199 4948 55255
rect 5004 55199 5014 55255
rect 4938 55113 4950 55199
rect 5002 55113 5014 55199
rect 4938 55057 4948 55113
rect 5004 55057 5014 55113
rect 4938 54971 4950 55057
rect 5002 54971 5014 55057
rect 4938 54915 4948 54971
rect 5004 54915 5014 54971
rect 4938 54829 4950 54915
rect 5002 54829 5014 54915
rect 4938 54773 4948 54829
rect 5004 54773 5014 54829
rect 4938 54687 4950 54773
rect 5002 54687 5014 54773
rect 4938 54631 4948 54687
rect 5004 54631 5014 54687
rect 4938 54624 4950 54631
rect 5002 54624 5014 54631
rect 4938 54612 5014 54624
rect 5426 55404 5502 55416
rect 5426 55397 5438 55404
rect 5490 55397 5502 55404
rect 5426 55341 5436 55397
rect 5492 55341 5502 55397
rect 5426 55255 5438 55341
rect 5490 55255 5502 55341
rect 5426 55199 5436 55255
rect 5492 55199 5502 55255
rect 5426 55113 5438 55199
rect 5490 55113 5502 55199
rect 5426 55057 5436 55113
rect 5492 55057 5502 55113
rect 5426 54971 5438 55057
rect 5490 54971 5502 55057
rect 5426 54915 5436 54971
rect 5492 54915 5502 54971
rect 5426 54829 5438 54915
rect 5490 54829 5502 54915
rect 5426 54773 5436 54829
rect 5492 54773 5502 54829
rect 5426 54687 5438 54773
rect 5490 54687 5502 54773
rect 5426 54631 5436 54687
rect 5492 54631 5502 54687
rect 5426 54624 5438 54631
rect 5490 54624 5502 54631
rect 5426 54612 5502 54624
rect 5914 55404 5990 55416
rect 5914 55397 5926 55404
rect 5978 55397 5990 55404
rect 5914 55341 5924 55397
rect 5980 55341 5990 55397
rect 6278 55404 6354 55416
rect 6278 55397 6290 55404
rect 6342 55397 6354 55404
rect 5914 55255 5926 55341
rect 5978 55255 5990 55341
rect 5914 55199 5924 55255
rect 5980 55199 5990 55255
rect 5914 55113 5926 55199
rect 5978 55113 5990 55199
rect 5914 55057 5924 55113
rect 5980 55057 5990 55113
rect 5914 54971 5926 55057
rect 5978 54971 5990 55057
rect 5914 54915 5924 54971
rect 5980 54915 5990 54971
rect 5914 54829 5926 54915
rect 5978 54829 5990 54915
rect 5914 54773 5924 54829
rect 5980 54773 5990 54829
rect 5914 54687 5926 54773
rect 5978 54687 5990 54773
rect 5914 54631 5924 54687
rect 5980 54631 5990 54687
rect 5914 54624 5926 54631
rect 5978 54624 5990 54631
rect 5914 54612 5990 54624
rect 6096 55371 6172 55381
rect 6096 55315 6106 55371
rect 6162 55315 6172 55371
rect 6096 55229 6108 55315
rect 6160 55229 6172 55315
rect 6096 55173 6106 55229
rect 6162 55173 6172 55229
rect 6096 55087 6108 55173
rect 6160 55087 6172 55173
rect 6096 55031 6106 55087
rect 6162 55031 6172 55087
rect 6096 54945 6108 55031
rect 6160 54945 6172 55031
rect 6096 54889 6106 54945
rect 6162 54889 6172 54945
rect 6096 54803 6108 54889
rect 6160 54803 6172 54889
rect 6096 54747 6106 54803
rect 6162 54747 6172 54803
rect 6096 54661 6108 54747
rect 6160 54661 6172 54747
rect 4162 54459 4238 54471
rect 6096 54605 6106 54661
rect 6162 54605 6172 54661
rect 6278 55341 6288 55397
rect 6344 55341 6354 55397
rect 6278 55255 6290 55341
rect 6342 55255 6354 55341
rect 6278 55199 6288 55255
rect 6344 55199 6354 55255
rect 6278 55113 6290 55199
rect 6342 55113 6354 55199
rect 6278 55057 6288 55113
rect 6344 55057 6354 55113
rect 6278 54971 6290 55057
rect 6342 54971 6354 55057
rect 6278 54915 6288 54971
rect 6344 54915 6354 54971
rect 6278 54829 6290 54915
rect 6342 54829 6354 54915
rect 6278 54773 6288 54829
rect 6344 54773 6354 54829
rect 6278 54687 6290 54773
rect 6342 54687 6354 54773
rect 6278 54631 6288 54687
rect 6344 54631 6354 54687
rect 6278 54624 6290 54631
rect 6342 54624 6354 54631
rect 6278 54612 6354 54624
rect 6766 55404 6842 55416
rect 6766 55397 6778 55404
rect 6830 55397 6842 55404
rect 6766 55341 6776 55397
rect 6832 55341 6842 55397
rect 6766 55255 6778 55341
rect 6830 55255 6842 55341
rect 6766 55199 6776 55255
rect 6832 55199 6842 55255
rect 6766 55113 6778 55199
rect 6830 55113 6842 55199
rect 6766 55057 6776 55113
rect 6832 55057 6842 55113
rect 6766 54971 6778 55057
rect 6830 54971 6842 55057
rect 6766 54915 6776 54971
rect 6832 54915 6842 54971
rect 6766 54829 6778 54915
rect 6830 54829 6842 54915
rect 6766 54773 6776 54829
rect 6832 54773 6842 54829
rect 6766 54687 6778 54773
rect 6830 54687 6842 54773
rect 6766 54631 6776 54687
rect 6832 54631 6842 54687
rect 6766 54624 6778 54631
rect 6830 54624 6842 54631
rect 6766 54612 6842 54624
rect 7254 55404 7330 55416
rect 7254 55397 7266 55404
rect 7318 55397 7330 55404
rect 7254 55341 7264 55397
rect 7320 55341 7330 55397
rect 7254 55255 7266 55341
rect 7318 55255 7330 55341
rect 7254 55199 7264 55255
rect 7320 55199 7330 55255
rect 7254 55113 7266 55199
rect 7318 55113 7330 55199
rect 7254 55057 7264 55113
rect 7320 55057 7330 55113
rect 7254 54971 7266 55057
rect 7318 54971 7330 55057
rect 7254 54915 7264 54971
rect 7320 54915 7330 54971
rect 7254 54829 7266 54915
rect 7318 54829 7330 54915
rect 7254 54773 7264 54829
rect 7320 54773 7330 54829
rect 7254 54687 7266 54773
rect 7318 54687 7330 54773
rect 7254 54631 7264 54687
rect 7320 54631 7330 54687
rect 7254 54624 7266 54631
rect 7318 54624 7330 54631
rect 7254 54612 7330 54624
rect 7434 55404 7510 55416
rect 7434 55397 7446 55404
rect 7498 55397 7510 55404
rect 7434 55341 7444 55397
rect 7500 55341 7510 55397
rect 7434 55255 7446 55341
rect 7498 55255 7510 55341
rect 7434 55199 7444 55255
rect 7500 55199 7510 55255
rect 7434 55113 7446 55199
rect 7498 55113 7510 55199
rect 7434 55057 7444 55113
rect 7500 55057 7510 55113
rect 7434 54971 7446 55057
rect 7498 54971 7510 55057
rect 7434 54915 7444 54971
rect 7500 54915 7510 54971
rect 7434 54829 7446 54915
rect 7498 54829 7510 54915
rect 7434 54773 7444 54829
rect 7500 54773 7510 54829
rect 7434 54687 7446 54773
rect 7498 54687 7510 54773
rect 7434 54631 7444 54687
rect 7500 54631 7510 54687
rect 7434 54624 7446 54631
rect 7498 54624 7510 54631
rect 7434 54612 7510 54624
rect 6096 54519 6108 54605
rect 6160 54519 6172 54605
rect 6096 54463 6106 54519
rect 6162 54463 6172 54519
rect 6096 54453 6172 54463
rect 8030 54471 8042 55459
rect 8094 54471 8106 55459
rect 8030 54459 8106 54471
rect 8499 55459 8575 55479
rect 8499 54471 8511 55459
rect 8563 54471 8575 55459
rect 8499 54459 8575 54471
rect 8714 55459 8790 55479
rect 8714 54471 8726 55459
rect 8778 54471 8790 55459
rect 8714 54459 8790 54471
rect 8937 55459 9013 55479
rect 8937 54471 8949 55459
rect 9001 54471 9013 55459
rect 8937 54459 9013 54471
rect 9406 55459 9482 55479
rect 9406 54471 9418 55459
rect 9470 54471 9482 55459
rect 13274 55459 13350 55479
rect 10002 55404 10078 55416
rect 10002 55397 10014 55404
rect 10066 55397 10078 55404
rect 10002 55341 10012 55397
rect 10068 55341 10078 55397
rect 10002 55255 10014 55341
rect 10066 55255 10078 55341
rect 10002 55199 10012 55255
rect 10068 55199 10078 55255
rect 10002 55113 10014 55199
rect 10066 55113 10078 55199
rect 10002 55057 10012 55113
rect 10068 55057 10078 55113
rect 10002 54971 10014 55057
rect 10066 54971 10078 55057
rect 10002 54915 10012 54971
rect 10068 54915 10078 54971
rect 10002 54829 10014 54915
rect 10066 54829 10078 54915
rect 10002 54773 10012 54829
rect 10068 54773 10078 54829
rect 10002 54687 10014 54773
rect 10066 54687 10078 54773
rect 10002 54631 10012 54687
rect 10068 54631 10078 54687
rect 10002 54624 10014 54631
rect 10066 54624 10078 54631
rect 10002 54612 10078 54624
rect 10182 55404 10258 55416
rect 10182 55397 10194 55404
rect 10246 55397 10258 55404
rect 10182 55341 10192 55397
rect 10248 55341 10258 55397
rect 10182 55255 10194 55341
rect 10246 55255 10258 55341
rect 10182 55199 10192 55255
rect 10248 55199 10258 55255
rect 10182 55113 10194 55199
rect 10246 55113 10258 55199
rect 10182 55057 10192 55113
rect 10248 55057 10258 55113
rect 10182 54971 10194 55057
rect 10246 54971 10258 55057
rect 10182 54915 10192 54971
rect 10248 54915 10258 54971
rect 10182 54829 10194 54915
rect 10246 54829 10258 54915
rect 10182 54773 10192 54829
rect 10248 54773 10258 54829
rect 10182 54687 10194 54773
rect 10246 54687 10258 54773
rect 10182 54631 10192 54687
rect 10248 54631 10258 54687
rect 10182 54624 10194 54631
rect 10246 54624 10258 54631
rect 10182 54612 10258 54624
rect 10670 55404 10746 55416
rect 10670 55397 10682 55404
rect 10734 55397 10746 55404
rect 10670 55341 10680 55397
rect 10736 55341 10746 55397
rect 10670 55255 10682 55341
rect 10734 55255 10746 55341
rect 10670 55199 10680 55255
rect 10736 55199 10746 55255
rect 10670 55113 10682 55199
rect 10734 55113 10746 55199
rect 10670 55057 10680 55113
rect 10736 55057 10746 55113
rect 10670 54971 10682 55057
rect 10734 54971 10746 55057
rect 10670 54915 10680 54971
rect 10736 54915 10746 54971
rect 10670 54829 10682 54915
rect 10734 54829 10746 54915
rect 10670 54773 10680 54829
rect 10736 54773 10746 54829
rect 10670 54687 10682 54773
rect 10734 54687 10746 54773
rect 10670 54631 10680 54687
rect 10736 54631 10746 54687
rect 10670 54624 10682 54631
rect 10734 54624 10746 54631
rect 10670 54612 10746 54624
rect 11158 55404 11234 55416
rect 11158 55397 11170 55404
rect 11222 55397 11234 55404
rect 11158 55341 11168 55397
rect 11224 55341 11234 55397
rect 11522 55404 11598 55416
rect 11522 55397 11534 55404
rect 11586 55397 11598 55404
rect 11158 55255 11170 55341
rect 11222 55255 11234 55341
rect 11158 55199 11168 55255
rect 11224 55199 11234 55255
rect 11158 55113 11170 55199
rect 11222 55113 11234 55199
rect 11158 55057 11168 55113
rect 11224 55057 11234 55113
rect 11158 54971 11170 55057
rect 11222 54971 11234 55057
rect 11158 54915 11168 54971
rect 11224 54915 11234 54971
rect 11158 54829 11170 54915
rect 11222 54829 11234 54915
rect 11158 54773 11168 54829
rect 11224 54773 11234 54829
rect 11158 54687 11170 54773
rect 11222 54687 11234 54773
rect 11158 54631 11168 54687
rect 11224 54631 11234 54687
rect 11158 54624 11170 54631
rect 11222 54624 11234 54631
rect 11158 54612 11234 54624
rect 11340 55371 11416 55381
rect 11340 55315 11350 55371
rect 11406 55315 11416 55371
rect 11340 55229 11352 55315
rect 11404 55229 11416 55315
rect 11340 55173 11350 55229
rect 11406 55173 11416 55229
rect 11340 55087 11352 55173
rect 11404 55087 11416 55173
rect 11340 55031 11350 55087
rect 11406 55031 11416 55087
rect 11340 54945 11352 55031
rect 11404 54945 11416 55031
rect 11340 54889 11350 54945
rect 11406 54889 11416 54945
rect 11340 54803 11352 54889
rect 11404 54803 11416 54889
rect 11340 54747 11350 54803
rect 11406 54747 11416 54803
rect 11340 54661 11352 54747
rect 11404 54661 11416 54747
rect 9406 54459 9482 54471
rect 11340 54605 11350 54661
rect 11406 54605 11416 54661
rect 11522 55341 11532 55397
rect 11588 55341 11598 55397
rect 11522 55255 11534 55341
rect 11586 55255 11598 55341
rect 11522 55199 11532 55255
rect 11588 55199 11598 55255
rect 11522 55113 11534 55199
rect 11586 55113 11598 55199
rect 11522 55057 11532 55113
rect 11588 55057 11598 55113
rect 11522 54971 11534 55057
rect 11586 54971 11598 55057
rect 11522 54915 11532 54971
rect 11588 54915 11598 54971
rect 11522 54829 11534 54915
rect 11586 54829 11598 54915
rect 11522 54773 11532 54829
rect 11588 54773 11598 54829
rect 11522 54687 11534 54773
rect 11586 54687 11598 54773
rect 11522 54631 11532 54687
rect 11588 54631 11598 54687
rect 11522 54624 11534 54631
rect 11586 54624 11598 54631
rect 11522 54612 11598 54624
rect 12010 55404 12086 55416
rect 12010 55397 12022 55404
rect 12074 55397 12086 55404
rect 12010 55341 12020 55397
rect 12076 55341 12086 55397
rect 12010 55255 12022 55341
rect 12074 55255 12086 55341
rect 12010 55199 12020 55255
rect 12076 55199 12086 55255
rect 12010 55113 12022 55199
rect 12074 55113 12086 55199
rect 12010 55057 12020 55113
rect 12076 55057 12086 55113
rect 12010 54971 12022 55057
rect 12074 54971 12086 55057
rect 12010 54915 12020 54971
rect 12076 54915 12086 54971
rect 12010 54829 12022 54915
rect 12074 54829 12086 54915
rect 12010 54773 12020 54829
rect 12076 54773 12086 54829
rect 12010 54687 12022 54773
rect 12074 54687 12086 54773
rect 12010 54631 12020 54687
rect 12076 54631 12086 54687
rect 12010 54624 12022 54631
rect 12074 54624 12086 54631
rect 12010 54612 12086 54624
rect 12498 55404 12574 55416
rect 12498 55397 12510 55404
rect 12562 55397 12574 55404
rect 12498 55341 12508 55397
rect 12564 55341 12574 55397
rect 12498 55255 12510 55341
rect 12562 55255 12574 55341
rect 12498 55199 12508 55255
rect 12564 55199 12574 55255
rect 12498 55113 12510 55199
rect 12562 55113 12574 55199
rect 12498 55057 12508 55113
rect 12564 55057 12574 55113
rect 12498 54971 12510 55057
rect 12562 54971 12574 55057
rect 12498 54915 12508 54971
rect 12564 54915 12574 54971
rect 12498 54829 12510 54915
rect 12562 54829 12574 54915
rect 12498 54773 12508 54829
rect 12564 54773 12574 54829
rect 12498 54687 12510 54773
rect 12562 54687 12574 54773
rect 12498 54631 12508 54687
rect 12564 54631 12574 54687
rect 12498 54624 12510 54631
rect 12562 54624 12574 54631
rect 12498 54612 12574 54624
rect 12678 55404 12754 55416
rect 12678 55397 12690 55404
rect 12742 55397 12754 55404
rect 12678 55341 12688 55397
rect 12744 55341 12754 55397
rect 12678 55255 12690 55341
rect 12742 55255 12754 55341
rect 12678 55199 12688 55255
rect 12744 55199 12754 55255
rect 12678 55113 12690 55199
rect 12742 55113 12754 55199
rect 12678 55057 12688 55113
rect 12744 55057 12754 55113
rect 12678 54971 12690 55057
rect 12742 54971 12754 55057
rect 12678 54915 12688 54971
rect 12744 54915 12754 54971
rect 12678 54829 12690 54915
rect 12742 54829 12754 54915
rect 12678 54773 12688 54829
rect 12744 54773 12754 54829
rect 12678 54687 12690 54773
rect 12742 54687 12754 54773
rect 12678 54631 12688 54687
rect 12744 54631 12754 54687
rect 12678 54624 12690 54631
rect 12742 54624 12754 54631
rect 12678 54612 12754 54624
rect 11340 54519 11352 54605
rect 11404 54519 11416 54605
rect 11340 54463 11350 54519
rect 11406 54463 11416 54519
rect 11340 54453 11416 54463
rect 13274 54471 13286 55459
rect 13338 54471 13350 55459
rect 13274 54459 13350 54471
rect 4162 54246 13350 54322
rect 3470 54001 3546 54013
rect 2098 53220 2347 53296
rect 1886 53087 1962 53173
rect 1886 53031 1896 53087
rect 1952 53031 1962 53087
rect 1886 52945 1962 53031
rect 1886 52889 1896 52945
rect 1952 52889 1962 52945
rect 1886 52803 1962 52889
rect 1886 52747 1896 52803
rect 1952 52747 1962 52803
rect 1886 52661 1962 52747
rect 1886 52605 1896 52661
rect 1952 52605 1962 52661
rect 3470 53013 3482 54001
rect 3534 53013 3546 54001
rect 4162 53793 4238 54246
rect 4162 53069 4174 53793
rect 3470 52649 3546 53013
rect 3788 53013 4174 53069
rect 4226 53013 4238 53793
rect 6096 53897 6172 53909
rect 6096 53814 6108 53897
rect 6160 53814 6172 53897
rect 6096 53758 6106 53814
rect 6162 53758 6172 53814
rect 3788 53001 4238 53013
rect 3788 52649 3895 53001
rect 4162 52999 4238 53001
rect 4758 53729 4834 53739
rect 4758 53673 4768 53729
rect 4824 53673 4834 53729
rect 4758 53632 4834 53673
rect 4758 53587 4770 53632
rect 4822 53587 4834 53632
rect 4758 53531 4768 53587
rect 4824 53531 4834 53587
rect 4758 53445 4770 53531
rect 4822 53445 4834 53531
rect 4758 53389 4768 53445
rect 4824 53389 4834 53445
rect 4758 53303 4770 53389
rect 4822 53303 4834 53389
rect 4758 53247 4768 53303
rect 4824 53247 4834 53303
rect 4758 53161 4770 53247
rect 4822 53161 4834 53247
rect 4758 53105 4768 53161
rect 4824 53105 4834 53161
rect 4758 53060 4770 53105
rect 4822 53060 4834 53105
rect 4758 53019 4834 53060
rect 4758 52963 4768 53019
rect 4824 52963 4834 53019
rect 4758 52953 4834 52963
rect 4938 53729 5014 53739
rect 4938 53673 4948 53729
rect 5004 53673 5014 53729
rect 4938 53632 5014 53673
rect 4938 53587 4950 53632
rect 5002 53587 5014 53632
rect 4938 53531 4948 53587
rect 5004 53531 5014 53587
rect 4938 53445 4950 53531
rect 5002 53445 5014 53531
rect 4938 53389 4948 53445
rect 5004 53389 5014 53445
rect 4938 53303 4950 53389
rect 5002 53303 5014 53389
rect 4938 53247 4948 53303
rect 5004 53247 5014 53303
rect 4938 53161 4950 53247
rect 5002 53161 5014 53247
rect 4938 53105 4948 53161
rect 5004 53105 5014 53161
rect 4938 53060 4950 53105
rect 5002 53060 5014 53105
rect 4938 53019 5014 53060
rect 4938 52963 4948 53019
rect 5004 52963 5014 53019
rect 4938 52953 5014 52963
rect 5426 53729 5502 53739
rect 5426 53673 5436 53729
rect 5492 53673 5502 53729
rect 5426 53632 5502 53673
rect 5426 53587 5438 53632
rect 5490 53587 5502 53632
rect 5426 53531 5436 53587
rect 5492 53531 5502 53587
rect 5426 53445 5438 53531
rect 5490 53445 5502 53531
rect 5426 53389 5436 53445
rect 5492 53389 5502 53445
rect 5426 53303 5438 53389
rect 5490 53303 5502 53389
rect 5426 53247 5436 53303
rect 5492 53247 5502 53303
rect 5426 53161 5438 53247
rect 5490 53161 5502 53247
rect 5426 53105 5436 53161
rect 5492 53105 5502 53161
rect 5426 53060 5438 53105
rect 5490 53060 5502 53105
rect 5426 53019 5502 53060
rect 5426 52963 5436 53019
rect 5492 52963 5502 53019
rect 5426 52953 5502 52963
rect 5914 53729 5990 53739
rect 5914 53673 5924 53729
rect 5980 53673 5990 53729
rect 5914 53632 5990 53673
rect 5914 53587 5926 53632
rect 5978 53587 5990 53632
rect 5914 53531 5924 53587
rect 5980 53531 5990 53587
rect 5914 53445 5926 53531
rect 5978 53445 5990 53531
rect 5914 53389 5924 53445
rect 5980 53389 5990 53445
rect 5914 53303 5926 53389
rect 5978 53303 5990 53389
rect 5914 53247 5924 53303
rect 5980 53247 5990 53303
rect 5914 53161 5926 53247
rect 5978 53161 5990 53247
rect 5914 53105 5924 53161
rect 5980 53105 5990 53161
rect 5914 53060 5926 53105
rect 5978 53060 5990 53105
rect 5914 53019 5990 53060
rect 5914 52963 5924 53019
rect 5980 52963 5990 53019
rect 5914 52953 5990 52963
rect 6096 53672 6108 53758
rect 6160 53672 6172 53758
rect 8030 53793 8106 54246
rect 6096 53616 6106 53672
rect 6162 53616 6172 53672
rect 6096 53530 6108 53616
rect 6160 53530 6172 53616
rect 6096 53474 6106 53530
rect 6162 53474 6172 53530
rect 6096 53388 6108 53474
rect 6160 53388 6172 53474
rect 6096 53332 6106 53388
rect 6162 53332 6172 53388
rect 6096 53246 6108 53332
rect 6160 53246 6172 53332
rect 6096 53190 6106 53246
rect 6162 53190 6172 53246
rect 6096 53104 6108 53190
rect 6160 53104 6172 53190
rect 6096 53048 6106 53104
rect 6162 53048 6172 53104
rect 6096 53013 6108 53048
rect 6160 53013 6172 53048
rect 6096 52962 6172 53013
rect 6096 52906 6106 52962
rect 6162 52906 6172 52962
rect 6278 53729 6354 53739
rect 6278 53673 6288 53729
rect 6344 53673 6354 53729
rect 6278 53632 6354 53673
rect 6278 53587 6290 53632
rect 6342 53587 6354 53632
rect 6278 53531 6288 53587
rect 6344 53531 6354 53587
rect 6278 53445 6290 53531
rect 6342 53445 6354 53531
rect 6278 53389 6288 53445
rect 6344 53389 6354 53445
rect 6278 53303 6290 53389
rect 6342 53303 6354 53389
rect 6278 53247 6288 53303
rect 6344 53247 6354 53303
rect 6278 53161 6290 53247
rect 6342 53161 6354 53247
rect 6278 53105 6288 53161
rect 6344 53105 6354 53161
rect 6278 53060 6290 53105
rect 6342 53060 6354 53105
rect 6278 53019 6354 53060
rect 6278 52963 6288 53019
rect 6344 52963 6354 53019
rect 6278 52953 6354 52963
rect 6766 53729 6842 53739
rect 6766 53673 6776 53729
rect 6832 53673 6842 53729
rect 6766 53632 6842 53673
rect 6766 53587 6778 53632
rect 6830 53587 6842 53632
rect 6766 53531 6776 53587
rect 6832 53531 6842 53587
rect 6766 53445 6778 53531
rect 6830 53445 6842 53531
rect 6766 53389 6776 53445
rect 6832 53389 6842 53445
rect 6766 53303 6778 53389
rect 6830 53303 6842 53389
rect 6766 53247 6776 53303
rect 6832 53247 6842 53303
rect 6766 53161 6778 53247
rect 6830 53161 6842 53247
rect 6766 53105 6776 53161
rect 6832 53105 6842 53161
rect 6766 53060 6778 53105
rect 6830 53060 6842 53105
rect 6766 53019 6842 53060
rect 6766 52963 6776 53019
rect 6832 52963 6842 53019
rect 6096 52896 6172 52906
rect 1886 52519 1962 52605
rect 3366 52637 3546 52649
rect 3366 52585 3378 52637
rect 3534 52585 3546 52637
rect 3366 52573 3546 52585
rect 3715 52637 3895 52649
rect 3715 52585 3727 52637
rect 3883 52585 3895 52637
rect 3715 52573 3895 52585
rect 1886 52463 1896 52519
rect 1952 52463 1962 52519
rect 1886 52453 1962 52463
rect 6766 52321 6842 52963
rect 7254 53729 7330 53739
rect 7254 53673 7264 53729
rect 7320 53673 7330 53729
rect 7254 53632 7330 53673
rect 7254 53587 7266 53632
rect 7318 53587 7330 53632
rect 7254 53531 7264 53587
rect 7320 53531 7330 53587
rect 7254 53445 7266 53531
rect 7318 53445 7330 53531
rect 7254 53389 7264 53445
rect 7320 53389 7330 53445
rect 7254 53303 7266 53389
rect 7318 53303 7330 53389
rect 7254 53247 7264 53303
rect 7320 53247 7330 53303
rect 7254 53161 7266 53247
rect 7318 53161 7330 53247
rect 7254 53105 7264 53161
rect 7320 53105 7330 53161
rect 7254 53060 7266 53105
rect 7318 53060 7330 53105
rect 7254 53019 7330 53060
rect 7254 52963 7264 53019
rect 7320 52963 7330 53019
rect 7254 52321 7330 52963
rect 7434 53729 7510 53739
rect 7434 53673 7444 53729
rect 7500 53673 7510 53729
rect 7434 53632 7510 53673
rect 7434 53587 7446 53632
rect 7498 53587 7510 53632
rect 7434 53531 7444 53587
rect 7500 53531 7510 53587
rect 7434 53445 7446 53531
rect 7498 53445 7510 53531
rect 7434 53389 7444 53445
rect 7500 53389 7510 53445
rect 7434 53303 7446 53389
rect 7498 53303 7510 53389
rect 7434 53247 7444 53303
rect 7500 53247 7510 53303
rect 7434 53161 7446 53247
rect 7498 53161 7510 53247
rect 7434 53105 7444 53161
rect 7500 53105 7510 53161
rect 7434 53060 7446 53105
rect 7498 53060 7510 53105
rect 7434 53019 7510 53060
rect 7434 52963 7444 53019
rect 7500 52963 7510 53019
rect 8030 53013 8042 53793
rect 8094 53013 8106 53793
rect 8030 53001 8106 53013
rect 8718 54001 8794 54246
rect 8718 53013 8730 54001
rect 8782 53013 8794 54001
rect 11340 53897 11416 53909
rect 7434 52953 7510 52963
rect 8718 52500 8794 53013
rect 9149 53797 9549 53830
rect 9149 53741 9179 53797
rect 9235 53741 9321 53797
rect 9377 53741 9463 53797
rect 9519 53741 9549 53797
rect 9149 53655 9549 53741
rect 11340 53814 11352 53897
rect 11404 53814 11416 53897
rect 11340 53758 11350 53814
rect 11406 53758 11416 53814
rect 9149 53599 9179 53655
rect 9235 53599 9321 53655
rect 9377 53599 9463 53655
rect 9519 53599 9549 53655
rect 9149 53513 9549 53599
rect 9149 53457 9179 53513
rect 9235 53457 9321 53513
rect 9377 53457 9463 53513
rect 9519 53457 9549 53513
rect 9149 53371 9549 53457
rect 9149 53315 9179 53371
rect 9235 53315 9321 53371
rect 9377 53315 9463 53371
rect 9519 53315 9549 53371
rect 9149 53229 9549 53315
rect 9149 53173 9179 53229
rect 9235 53173 9321 53229
rect 9377 53173 9463 53229
rect 9519 53173 9549 53229
rect 9149 53087 9549 53173
rect 9149 53031 9179 53087
rect 9235 53031 9321 53087
rect 9377 53031 9463 53087
rect 9519 53031 9549 53087
rect 9149 52945 9549 53031
rect 10002 53729 10078 53739
rect 10002 53673 10012 53729
rect 10068 53673 10078 53729
rect 10002 53632 10078 53673
rect 10002 53587 10014 53632
rect 10066 53587 10078 53632
rect 10002 53531 10012 53587
rect 10068 53531 10078 53587
rect 10002 53445 10014 53531
rect 10066 53445 10078 53531
rect 10002 53389 10012 53445
rect 10068 53389 10078 53445
rect 10002 53303 10014 53389
rect 10066 53303 10078 53389
rect 10002 53247 10012 53303
rect 10068 53247 10078 53303
rect 10002 53161 10014 53247
rect 10066 53161 10078 53247
rect 10002 53105 10012 53161
rect 10068 53105 10078 53161
rect 10002 53060 10014 53105
rect 10066 53060 10078 53105
rect 10002 53019 10078 53060
rect 10002 52963 10012 53019
rect 10068 52963 10078 53019
rect 10002 52953 10078 52963
rect 10182 53729 10258 53739
rect 10182 53673 10192 53729
rect 10248 53673 10258 53729
rect 10182 53632 10258 53673
rect 10182 53587 10194 53632
rect 10246 53587 10258 53632
rect 10182 53531 10192 53587
rect 10248 53531 10258 53587
rect 10182 53445 10194 53531
rect 10246 53445 10258 53531
rect 10182 53389 10192 53445
rect 10248 53389 10258 53445
rect 10182 53303 10194 53389
rect 10246 53303 10258 53389
rect 10182 53247 10192 53303
rect 10248 53247 10258 53303
rect 10182 53161 10194 53247
rect 10246 53161 10258 53247
rect 10182 53105 10192 53161
rect 10248 53105 10258 53161
rect 10182 53060 10194 53105
rect 10246 53060 10258 53105
rect 10182 53019 10258 53060
rect 10182 52963 10192 53019
rect 10248 52963 10258 53019
rect 10182 52953 10258 52963
rect 10670 53729 10746 53739
rect 10670 53673 10680 53729
rect 10736 53673 10746 53729
rect 10670 53632 10746 53673
rect 10670 53587 10682 53632
rect 10734 53587 10746 53632
rect 10670 53531 10680 53587
rect 10736 53531 10746 53587
rect 10670 53445 10682 53531
rect 10734 53445 10746 53531
rect 10670 53389 10680 53445
rect 10736 53389 10746 53445
rect 10670 53303 10682 53389
rect 10734 53303 10746 53389
rect 10670 53247 10680 53303
rect 10736 53247 10746 53303
rect 10670 53161 10682 53247
rect 10734 53161 10746 53247
rect 10670 53105 10680 53161
rect 10736 53105 10746 53161
rect 10670 53060 10682 53105
rect 10734 53060 10746 53105
rect 10670 53019 10746 53060
rect 10670 52963 10680 53019
rect 10736 52963 10746 53019
rect 10670 52953 10746 52963
rect 11158 53729 11234 53739
rect 11158 53673 11168 53729
rect 11224 53673 11234 53729
rect 11158 53632 11234 53673
rect 11158 53587 11170 53632
rect 11222 53587 11234 53632
rect 11158 53531 11168 53587
rect 11224 53531 11234 53587
rect 11158 53445 11170 53531
rect 11222 53445 11234 53531
rect 11158 53389 11168 53445
rect 11224 53389 11234 53445
rect 11158 53303 11170 53389
rect 11222 53303 11234 53389
rect 11158 53247 11168 53303
rect 11224 53247 11234 53303
rect 11158 53161 11170 53247
rect 11222 53161 11234 53247
rect 11158 53105 11168 53161
rect 11224 53105 11234 53161
rect 11158 53060 11170 53105
rect 11222 53060 11234 53105
rect 11158 53019 11234 53060
rect 11158 52963 11168 53019
rect 11224 52963 11234 53019
rect 11158 52953 11234 52963
rect 11340 53672 11352 53758
rect 11404 53672 11416 53758
rect 13274 53793 13350 54246
rect 11340 53616 11350 53672
rect 11406 53616 11416 53672
rect 11340 53530 11352 53616
rect 11404 53530 11416 53616
rect 11340 53474 11350 53530
rect 11406 53474 11416 53530
rect 11340 53388 11352 53474
rect 11404 53388 11416 53474
rect 11340 53332 11350 53388
rect 11406 53332 11416 53388
rect 11340 53246 11352 53332
rect 11404 53246 11416 53332
rect 11340 53190 11350 53246
rect 11406 53190 11416 53246
rect 11340 53104 11352 53190
rect 11404 53104 11416 53190
rect 11340 53048 11350 53104
rect 11406 53048 11416 53104
rect 11340 53013 11352 53048
rect 11404 53013 11416 53048
rect 11340 52962 11416 53013
rect 9149 52889 9179 52945
rect 9235 52889 9321 52945
rect 9377 52889 9463 52945
rect 9519 52889 9549 52945
rect 11340 52906 11350 52962
rect 11406 52906 11416 52962
rect 11522 53729 11598 53739
rect 11522 53673 11532 53729
rect 11588 53673 11598 53729
rect 11522 53632 11598 53673
rect 11522 53587 11534 53632
rect 11586 53587 11598 53632
rect 11522 53531 11532 53587
rect 11588 53531 11598 53587
rect 11522 53445 11534 53531
rect 11586 53445 11598 53531
rect 11522 53389 11532 53445
rect 11588 53389 11598 53445
rect 11522 53303 11534 53389
rect 11586 53303 11598 53389
rect 11522 53247 11532 53303
rect 11588 53247 11598 53303
rect 11522 53161 11534 53247
rect 11586 53161 11598 53247
rect 11522 53105 11532 53161
rect 11588 53105 11598 53161
rect 11522 53060 11534 53105
rect 11586 53060 11598 53105
rect 11522 53019 11598 53060
rect 11522 52963 11532 53019
rect 11588 52963 11598 53019
rect 11522 52953 11598 52963
rect 12010 53729 12086 53739
rect 12010 53673 12020 53729
rect 12076 53673 12086 53729
rect 12010 53632 12086 53673
rect 12010 53587 12022 53632
rect 12074 53587 12086 53632
rect 12010 53531 12020 53587
rect 12076 53531 12086 53587
rect 12010 53445 12022 53531
rect 12074 53445 12086 53531
rect 12010 53389 12020 53445
rect 12076 53389 12086 53445
rect 12010 53303 12022 53389
rect 12074 53303 12086 53389
rect 12010 53247 12020 53303
rect 12076 53247 12086 53303
rect 12010 53161 12022 53247
rect 12074 53161 12086 53247
rect 12010 53105 12020 53161
rect 12076 53105 12086 53161
rect 12010 53060 12022 53105
rect 12074 53060 12086 53105
rect 12010 53019 12086 53060
rect 12010 52963 12020 53019
rect 12076 52963 12086 53019
rect 12010 52953 12086 52963
rect 12498 53729 12574 53739
rect 12498 53673 12508 53729
rect 12564 53673 12574 53729
rect 12498 53632 12574 53673
rect 12498 53587 12510 53632
rect 12562 53587 12574 53632
rect 12498 53531 12508 53587
rect 12564 53531 12574 53587
rect 12498 53445 12510 53531
rect 12562 53445 12574 53531
rect 12498 53389 12508 53445
rect 12564 53389 12574 53445
rect 12498 53303 12510 53389
rect 12562 53303 12574 53389
rect 12498 53247 12508 53303
rect 12564 53247 12574 53303
rect 12498 53161 12510 53247
rect 12562 53161 12574 53247
rect 12498 53105 12508 53161
rect 12564 53105 12574 53161
rect 12498 53060 12510 53105
rect 12562 53060 12574 53105
rect 12498 53019 12574 53060
rect 12498 52963 12508 53019
rect 12564 52963 12574 53019
rect 12498 52953 12574 52963
rect 12678 53729 12754 53739
rect 12678 53673 12688 53729
rect 12744 53673 12754 53729
rect 12678 53632 12754 53673
rect 12678 53587 12690 53632
rect 12742 53587 12754 53632
rect 12678 53531 12688 53587
rect 12744 53531 12754 53587
rect 12678 53445 12690 53531
rect 12742 53445 12754 53531
rect 12678 53389 12688 53445
rect 12744 53389 12754 53445
rect 12678 53303 12690 53389
rect 12742 53303 12754 53389
rect 12678 53247 12688 53303
rect 12744 53247 12754 53303
rect 12678 53161 12690 53247
rect 12742 53161 12754 53247
rect 12678 53105 12688 53161
rect 12744 53105 12754 53161
rect 12678 53060 12690 53105
rect 12742 53060 12754 53105
rect 12678 53019 12754 53060
rect 12678 52963 12688 53019
rect 12744 52963 12754 53019
rect 13274 53013 13286 53793
rect 13338 53013 13350 53793
rect 13274 53001 13350 53013
rect 12678 52953 12754 52963
rect 11340 52896 11416 52906
rect 9149 52803 9549 52889
rect 9149 52747 9179 52803
rect 9235 52747 9321 52803
rect 9377 52747 9463 52803
rect 9519 52747 9549 52803
rect 9149 52661 9549 52747
rect 9149 52605 9179 52661
rect 9235 52605 9321 52661
rect 9377 52605 9463 52661
rect 9519 52605 9549 52661
rect 9149 52519 9549 52605
rect 9149 52463 9179 52519
rect 9235 52463 9321 52519
rect 9377 52463 9463 52519
rect 9519 52463 9549 52519
rect 9149 52407 9549 52463
rect 6438 52309 6930 52321
rect 6438 52257 6450 52309
rect 6918 52257 6930 52309
rect 6438 52245 6930 52257
rect 7254 52309 9010 52321
rect 7254 52257 7266 52309
rect 7422 52257 9010 52309
rect 7254 52237 9010 52257
rect 9149 50960 9428 52407
rect 2528 49899 6140 49911
rect 2528 49847 2540 49899
rect 6128 49847 6140 49899
rect 2528 49835 6140 49847
rect 7714 49899 8114 49911
rect 7714 49847 7732 49899
rect 8096 49847 8114 49899
rect 4594 49054 4994 49835
rect 4594 49002 4644 49054
rect 4696 49002 4768 49054
rect 4820 49002 4892 49054
rect 4944 49002 4994 49054
rect 4594 48930 4994 49002
rect 3978 48918 4302 48928
rect 3978 48862 3988 48918
rect 4044 48862 4112 48918
rect 4168 48862 4236 48918
rect 4292 48862 4302 48918
rect 3978 48794 4302 48862
rect 3978 48738 3988 48794
rect 4044 48738 4112 48794
rect 4168 48738 4236 48794
rect 4292 48738 4302 48794
rect 3978 48670 4302 48738
rect 3978 48614 3988 48670
rect 4044 48614 4112 48670
rect 4168 48614 4236 48670
rect 4292 48614 4302 48670
rect 3978 48546 4302 48614
rect 3978 48490 3988 48546
rect 4044 48490 4112 48546
rect 4168 48490 4236 48546
rect 4292 48490 4302 48546
rect 3978 48422 4302 48490
rect 3978 48366 3988 48422
rect 4044 48366 4112 48422
rect 4168 48366 4236 48422
rect 4292 48366 4302 48422
rect 3978 48298 4302 48366
rect 3978 48242 3988 48298
rect 4044 48242 4112 48298
rect 4168 48242 4236 48298
rect 4292 48242 4302 48298
rect 3978 48174 4302 48242
rect 3978 48118 3988 48174
rect 4044 48118 4112 48174
rect 4168 48118 4236 48174
rect 4292 48118 4302 48174
rect 3978 48050 4302 48118
rect 3978 47994 3988 48050
rect 4044 47994 4112 48050
rect 4168 47994 4236 48050
rect 4292 47994 4302 48050
rect 3978 47926 4302 47994
rect 3978 47870 3988 47926
rect 4044 47870 4112 47926
rect 4168 47870 4236 47926
rect 4292 47870 4302 47926
rect 3978 47802 4302 47870
rect 3978 47746 3988 47802
rect 4044 47746 4112 47802
rect 4168 47746 4236 47802
rect 4292 47746 4302 47802
rect 3978 47736 4302 47746
rect 4594 48878 4644 48930
rect 4696 48878 4768 48930
rect 4820 48878 4892 48930
rect 4944 48878 4994 48930
rect 4594 48806 4994 48878
rect 4594 48754 4644 48806
rect 4696 48754 4768 48806
rect 4820 48754 4892 48806
rect 4944 48754 4994 48806
rect 4594 48682 4994 48754
rect 5513 49028 5913 49835
rect 5513 48768 5531 49028
rect 5895 48768 5913 49028
rect 5513 48710 5913 48768
rect 4594 48630 4644 48682
rect 4696 48630 4768 48682
rect 4820 48630 4892 48682
rect 4944 48630 4994 48682
rect 4594 48558 4994 48630
rect 4594 48506 4644 48558
rect 4696 48506 4768 48558
rect 4820 48506 4892 48558
rect 4944 48506 4994 48558
rect 4594 48434 4994 48506
rect 4594 48382 4644 48434
rect 4696 48382 4768 48434
rect 4820 48382 4892 48434
rect 4944 48382 4994 48434
rect 4594 48310 4994 48382
rect 4594 48258 4644 48310
rect 4696 48258 4768 48310
rect 4820 48258 4892 48310
rect 4944 48258 4994 48310
rect 4594 48186 4994 48258
rect 4594 48134 4644 48186
rect 4696 48134 4768 48186
rect 4820 48134 4892 48186
rect 4944 48134 4994 48186
rect 4594 48062 4994 48134
rect 4594 48010 4644 48062
rect 4696 48010 4768 48062
rect 4820 48010 4892 48062
rect 4944 48010 4994 48062
rect 4594 47938 4994 48010
rect 4594 47886 4644 47938
rect 4696 47886 4768 47938
rect 4820 47886 4892 47938
rect 4944 47886 4994 47938
rect 4594 47814 4994 47886
rect 4594 47762 4644 47814
rect 4696 47762 4768 47814
rect 4820 47762 4892 47814
rect 4944 47762 4994 47814
rect 4594 47690 4994 47762
rect 4594 47638 4644 47690
rect 4696 47638 4768 47690
rect 4820 47638 4892 47690
rect 4944 47638 4994 47690
rect 4594 47566 4994 47638
rect 4594 47514 4644 47566
rect 4696 47514 4768 47566
rect 4820 47514 4892 47566
rect 4944 47514 4994 47566
rect 3608 47418 3684 47430
rect 3608 47414 3620 47418
rect 3672 47414 3684 47418
rect 3608 47358 3618 47414
rect 3674 47358 3684 47414
rect 3608 47272 3620 47358
rect 3672 47272 3684 47358
rect 3608 47216 3618 47272
rect 3674 47216 3684 47272
rect 3608 47130 3620 47216
rect 3672 47130 3684 47216
rect 3608 47074 3618 47130
rect 3674 47074 3684 47130
rect 3608 46988 3620 47074
rect 3672 46988 3684 47074
rect 3608 46932 3618 46988
rect 3674 46932 3684 46988
rect 3608 46846 3620 46932
rect 3672 46846 3684 46932
rect 3608 46790 3618 46846
rect 3674 46790 3684 46846
rect 3608 46704 3620 46790
rect 3672 46704 3684 46790
rect 3608 46648 3618 46704
rect 3674 46648 3684 46704
rect 3608 46562 3620 46648
rect 3672 46562 3684 46648
rect 3608 46506 3618 46562
rect 3674 46506 3684 46562
rect 3608 46420 3620 46506
rect 3672 46420 3684 46506
rect 3608 46364 3618 46420
rect 3674 46364 3684 46420
rect 3608 46326 3620 46364
rect 3672 46326 3684 46364
rect 3608 46314 3684 46326
rect 4594 46250 4994 47514
rect 3158 46134 4378 46150
rect 3158 45666 3197 46134
rect 3353 45666 4378 46134
rect 3158 45650 4378 45666
rect 7427 45650 7627 49191
rect 7714 49028 8114 49847
rect 7714 48768 7732 49028
rect 8096 48768 8114 49028
rect 7714 48710 8114 48768
rect 8416 49899 8816 49911
rect 8416 49847 8434 49899
rect 8798 49847 8816 49899
rect 8416 49028 8816 49847
rect 8416 48768 8434 49028
rect 8798 48768 8816 49028
rect 8416 48710 8816 48768
rect 9149 48292 9549 50960
rect 11552 49568 11740 49578
rect 11552 49512 11562 49568
rect 11618 49512 11674 49568
rect 11730 49512 11740 49568
rect 11552 49456 11740 49512
rect 11552 49400 11562 49456
rect 11618 49400 11674 49456
rect 11730 49400 11740 49456
rect 11552 49344 11740 49400
rect 11552 49288 11562 49344
rect 11618 49288 11674 49344
rect 11730 49288 11740 49344
rect 11552 49278 11740 49288
rect 10782 49014 10858 49024
rect 10782 48958 10792 49014
rect 10848 48958 10858 49014
rect 10782 48872 10794 48958
rect 10846 48872 10858 48958
rect 10782 48816 10792 48872
rect 10848 48816 10858 48872
rect 10782 48730 10794 48816
rect 10846 48730 10858 48816
rect 10782 48674 10792 48730
rect 10848 48674 10858 48730
rect 10782 48588 10794 48674
rect 10846 48588 10858 48674
rect 10782 48532 10792 48588
rect 10848 48532 10858 48588
rect 10782 48446 10794 48532
rect 10846 48446 10858 48532
rect 10782 48390 10792 48446
rect 10848 48390 10858 48446
rect 10782 48304 10794 48390
rect 10846 48304 10858 48390
rect 10782 48248 10792 48304
rect 10848 48248 10858 48304
rect 10782 48162 10794 48248
rect 10846 48162 10858 48248
rect 10782 48106 10792 48162
rect 10848 48106 10858 48162
rect 10782 48020 10794 48106
rect 10846 48020 10858 48106
rect 10782 47964 10792 48020
rect 10848 47964 10858 48020
rect 10782 47954 10858 47964
rect 9713 45830 9931 47661
rect 11567 47608 11720 49278
rect 11567 47452 11608 47608
rect 11660 47452 11720 47608
rect 11567 47440 11720 47452
rect 11001 47404 11077 47416
rect 11001 47397 11013 47404
rect 11065 47397 11077 47404
rect 11001 47341 11011 47397
rect 11067 47341 11077 47397
rect 11001 47255 11013 47341
rect 11065 47255 11077 47341
rect 11001 47199 11011 47255
rect 11067 47199 11077 47255
rect 11001 47113 11013 47199
rect 11065 47113 11077 47199
rect 11001 47057 11011 47113
rect 11067 47057 11077 47113
rect 11001 46971 11013 47057
rect 11065 46971 11077 47057
rect 11001 46915 11011 46971
rect 11067 46915 11077 46971
rect 11001 46829 11013 46915
rect 11065 46829 11077 46915
rect 11001 46773 11011 46829
rect 11067 46773 11077 46829
rect 11001 46687 11013 46773
rect 11065 46687 11077 46773
rect 11001 46631 11011 46687
rect 11067 46631 11077 46687
rect 11001 46624 11013 46631
rect 11065 46624 11077 46631
rect 11001 46612 11077 46624
rect 3969 45341 4293 45351
rect 3969 45285 3979 45341
rect 4035 45285 4103 45341
rect 4159 45285 4227 45341
rect 4283 45285 4293 45341
rect 3969 45217 4293 45285
rect 3969 45161 3979 45217
rect 4035 45161 4103 45217
rect 4159 45161 4227 45217
rect 4283 45161 4293 45217
rect 3969 45093 4293 45161
rect 3969 45037 3979 45093
rect 4035 45037 4103 45093
rect 4159 45037 4227 45093
rect 4283 45037 4293 45093
rect 3969 44969 4293 45037
rect 3969 44913 3979 44969
rect 4035 44913 4103 44969
rect 4159 44913 4227 44969
rect 4283 44913 4293 44969
rect 3969 44845 4293 44913
rect 3969 44789 3979 44845
rect 4035 44789 4103 44845
rect 4159 44789 4227 44845
rect 4283 44789 4293 44845
rect 3969 44721 4293 44789
rect 3969 44665 3979 44721
rect 4035 44665 4103 44721
rect 4159 44665 4227 44721
rect 4283 44665 4293 44721
rect 3969 44597 4293 44665
rect 3969 44541 3979 44597
rect 4035 44541 4103 44597
rect 4159 44541 4227 44597
rect 4283 44541 4293 44597
rect 3969 44531 4293 44541
rect 9713 44430 10470 45830
rect 3608 44197 3684 44207
rect 3608 44141 3618 44197
rect 3674 44141 3684 44197
rect 3608 44055 3620 44141
rect 3672 44055 3684 44141
rect 3608 43999 3618 44055
rect 3674 43999 3684 44055
rect 3608 43913 3620 43999
rect 3672 43913 3684 43999
rect 3608 43857 3618 43913
rect 3674 43857 3684 43913
rect 3608 43771 3620 43857
rect 3672 43771 3684 43857
rect 3608 43715 3618 43771
rect 3674 43715 3684 43771
rect 3608 43629 3620 43715
rect 3672 43629 3684 43715
rect 3608 43573 3618 43629
rect 3674 43573 3684 43629
rect 3608 43487 3620 43573
rect 3672 43487 3684 43573
rect 3608 43431 3618 43487
rect 3674 43431 3684 43487
rect 3608 43345 3620 43431
rect 3672 43345 3684 43431
rect 3608 43289 3618 43345
rect 3674 43289 3684 43345
rect 3608 43203 3620 43289
rect 3672 43203 3684 43289
rect 3608 43147 3618 43203
rect 3674 43147 3684 43203
rect 3608 43061 3620 43147
rect 3672 43061 3684 43147
rect 3608 43005 3618 43061
rect 3674 43005 3684 43061
rect 3608 42919 3620 43005
rect 3672 42919 3684 43005
rect 3608 42863 3618 42919
rect 3674 42863 3684 42919
rect 3608 42853 3684 42863
rect 12406 43683 12624 43695
rect 12406 43631 12437 43683
rect 12593 43631 12624 43683
rect 3608 42597 3684 42607
rect 3608 42541 3618 42597
rect 3674 42541 3684 42597
rect 3608 42455 3620 42541
rect 3672 42455 3684 42541
rect 3608 42399 3618 42455
rect 3674 42399 3684 42455
rect 3608 42313 3620 42399
rect 3672 42313 3684 42399
rect 3608 42257 3618 42313
rect 3674 42257 3684 42313
rect 3608 42171 3620 42257
rect 3672 42171 3684 42257
rect 3608 42115 3618 42171
rect 3674 42115 3684 42171
rect 3608 42029 3620 42115
rect 3672 42029 3684 42115
rect 3608 41973 3618 42029
rect 3674 41973 3684 42029
rect 3608 41887 3620 41973
rect 3672 41887 3684 41973
rect 3608 41831 3618 41887
rect 3674 41831 3684 41887
rect 3608 41745 3620 41831
rect 3672 41745 3684 41831
rect 3608 41689 3618 41745
rect 3674 41689 3684 41745
rect 3608 41603 3620 41689
rect 3672 41603 3684 41689
rect 3608 41547 3618 41603
rect 3674 41547 3684 41603
rect 3608 41461 3620 41547
rect 3672 41461 3684 41547
rect 3608 41405 3618 41461
rect 3674 41405 3684 41461
rect 3608 41319 3620 41405
rect 3672 41319 3684 41405
rect 3608 41263 3618 41319
rect 3674 41263 3684 41319
rect 11356 41444 11581 41456
rect 3608 41253 3684 41263
rect 1836 40702 3758 40712
rect 1836 40646 1846 40702
rect 1902 40700 1988 40702
rect 2044 40700 2130 40702
rect 2186 40700 2272 40702
rect 2328 40700 2414 40702
rect 2470 40700 2556 40702
rect 2612 40700 2698 40702
rect 2754 40700 2840 40702
rect 2896 40700 2982 40702
rect 3038 40700 3124 40702
rect 3180 40700 3266 40702
rect 3322 40700 3408 40702
rect 3464 40700 3550 40702
rect 3606 40700 3692 40702
rect 3668 40648 3692 40700
rect 1902 40646 1988 40648
rect 2044 40646 2130 40648
rect 2186 40646 2272 40648
rect 2328 40646 2414 40648
rect 2470 40646 2556 40648
rect 2612 40646 2698 40648
rect 2754 40646 2840 40648
rect 2896 40646 2982 40648
rect 3038 40646 3124 40648
rect 3180 40646 3266 40648
rect 3322 40646 3408 40648
rect 3464 40646 3550 40648
rect 3606 40646 3692 40648
rect 3748 40646 3758 40702
rect 1836 40636 3758 40646
rect 1913 40364 2093 40376
rect 1913 40312 1925 40364
rect 2081 40312 2093 40364
rect 1913 40300 2093 40312
rect 4837 40364 5017 40376
rect 4837 40312 4849 40364
rect 5005 40312 5017 40364
rect 4837 40300 5017 40312
rect 7053 40364 7233 40376
rect 7053 40312 7065 40364
rect 7221 40312 7233 40364
rect 7053 40300 7233 40312
rect 1596 40228 1776 40240
rect 1596 40176 1608 40228
rect 1764 40176 1776 40228
rect 1596 40164 1776 40176
rect 1184 38687 1260 40163
rect 1771 39420 1847 39430
rect 1771 39364 1781 39420
rect 1837 39364 1847 39420
rect 1771 39278 1783 39364
rect 1835 39278 1847 39364
rect 1771 39222 1781 39278
rect 1837 39222 1847 39278
rect 1771 39136 1783 39222
rect 1835 39136 1847 39222
rect 1771 39080 1781 39136
rect 1837 39080 1847 39136
rect 1771 38994 1783 39080
rect 1835 38994 1847 39080
rect 1771 38938 1781 38994
rect 1837 38938 1847 38994
rect 1771 38852 1783 38938
rect 1835 38852 1847 38938
rect 1771 38796 1781 38852
rect 1837 38796 1847 38852
rect 1771 38786 1847 38796
rect 1913 38687 1989 40300
rect 2428 39946 4492 39956
rect 2428 39890 2438 39946
rect 2494 39944 2580 39946
rect 2636 39944 2722 39946
rect 2778 39944 2864 39946
rect 2920 39944 3006 39946
rect 3062 39944 3148 39946
rect 3204 39944 3290 39946
rect 3346 39944 3432 39946
rect 3488 39944 3574 39946
rect 3630 39944 3716 39946
rect 3772 39944 3858 39946
rect 3914 39944 4000 39946
rect 4056 39944 4142 39946
rect 4198 39944 4284 39946
rect 4340 39944 4426 39946
rect 2494 39890 2580 39892
rect 2636 39890 2722 39892
rect 2778 39890 2864 39892
rect 2920 39890 3006 39892
rect 3062 39890 3148 39892
rect 3204 39890 3290 39892
rect 3346 39890 3432 39892
rect 3488 39890 3574 39892
rect 3630 39890 3716 39892
rect 3772 39890 3858 39892
rect 3914 39890 4000 39892
rect 4056 39890 4142 39892
rect 4198 39890 4284 39892
rect 4340 39890 4426 39892
rect 4482 39890 4492 39946
rect 2428 39880 4492 39890
rect 4941 38687 5017 40300
rect 5566 40228 5746 40240
rect 5566 40176 5578 40228
rect 5734 40176 5746 40228
rect 5566 40164 5746 40176
rect 5083 39420 5159 39430
rect 5083 39364 5093 39420
rect 5149 39364 5159 39420
rect 5083 39278 5095 39364
rect 5147 39278 5159 39364
rect 5083 39222 5093 39278
rect 5149 39222 5159 39278
rect 5083 39136 5095 39222
rect 5147 39136 5159 39222
rect 5083 39080 5093 39136
rect 5149 39080 5159 39136
rect 5083 38994 5095 39080
rect 5147 38994 5159 39080
rect 5083 38938 5093 38994
rect 5149 38938 5159 38994
rect 5083 38852 5095 38938
rect 5147 38852 5159 38938
rect 5083 38796 5093 38852
rect 5149 38796 5159 38852
rect 5083 38786 5159 38796
rect 5670 38687 5746 40164
rect 6049 39418 6125 39430
rect 6049 39414 6061 39418
rect 6113 39414 6125 39418
rect 6049 39358 6059 39414
rect 6115 39358 6125 39414
rect 6049 39272 6061 39358
rect 6113 39272 6125 39358
rect 6049 39216 6059 39272
rect 6115 39216 6125 39272
rect 6049 39130 6061 39216
rect 6113 39130 6125 39216
rect 6049 39074 6059 39130
rect 6115 39074 6125 39130
rect 6049 38988 6061 39074
rect 6113 38988 6125 39074
rect 6049 38932 6059 38988
rect 6115 38932 6125 38988
rect 6049 38846 6061 38932
rect 6113 38846 6125 38932
rect 6049 38790 6059 38846
rect 6115 38790 6125 38846
rect 6049 38704 6061 38790
rect 6113 38704 6125 38790
rect 7015 39420 7091 39430
rect 7015 39364 7025 39420
rect 7081 39364 7091 39420
rect 7015 39278 7027 39364
rect 7079 39278 7091 39364
rect 7015 39222 7025 39278
rect 7081 39222 7091 39278
rect 7015 39136 7027 39222
rect 7079 39136 7091 39222
rect 7015 39080 7025 39136
rect 7081 39080 7091 39136
rect 7015 38994 7027 39080
rect 7079 38994 7091 39080
rect 7015 38938 7025 38994
rect 7081 38938 7091 38994
rect 7015 38852 7027 38938
rect 7079 38852 7091 38938
rect 7015 38796 7025 38852
rect 7081 38796 7091 38852
rect 7015 38786 7091 38796
rect 6049 38648 6059 38704
rect 6115 38648 6125 38704
rect 7157 38687 7233 40300
rect 6049 38562 6061 38648
rect 6113 38562 6125 38648
rect 6049 38506 6059 38562
rect 6115 38506 6125 38562
rect 6049 38430 6061 38506
rect 6113 38430 6125 38506
rect 6049 38420 6125 38430
rect 6049 38364 6059 38420
rect 6115 38364 6125 38420
rect 6049 38354 6125 38364
rect 32 37797 122 37830
rect 32 37741 56 37797
rect 112 37741 122 37797
rect 32 37655 58 37741
rect 110 37655 122 37741
rect 32 37599 56 37655
rect 112 37599 122 37655
rect 32 37513 58 37599
rect 110 37513 122 37599
rect 32 37457 56 37513
rect 112 37457 122 37513
rect 32 37371 58 37457
rect 110 37371 122 37457
rect 32 37315 56 37371
rect 112 37315 122 37371
rect 32 37229 58 37315
rect 110 37229 122 37315
rect 32 37173 56 37229
rect 112 37173 122 37229
rect 32 37087 58 37173
rect 110 37087 122 37173
rect 32 37031 56 37087
rect 112 37031 122 37087
rect 32 36945 58 37031
rect 110 36945 122 37031
rect 32 36889 56 36945
rect 112 36889 122 36945
rect 32 36803 58 36889
rect 110 36803 122 36889
rect 32 36747 56 36803
rect 112 36747 122 36803
rect 32 36661 58 36747
rect 110 36661 122 36747
rect 32 36605 56 36661
rect 112 36605 122 36661
rect 32 36519 58 36605
rect 110 36519 122 36605
rect 32 36463 56 36519
rect 112 36463 122 36519
rect 32 36430 122 36463
rect 704 37797 817 38142
rect 704 37741 734 37797
rect 790 37741 817 37797
rect 704 37655 817 37741
rect 704 37599 734 37655
rect 790 37599 817 37655
rect 704 37513 817 37599
rect 704 37457 734 37513
rect 790 37457 817 37513
rect 704 37371 817 37457
rect 704 37315 734 37371
rect 790 37315 817 37371
rect 704 37229 817 37315
rect 704 37173 734 37229
rect 790 37173 817 37229
rect 704 37154 817 37173
rect 869 37797 1104 38142
rect 869 37741 876 37797
rect 932 37741 1018 37797
rect 1074 37741 1104 37797
rect 869 37655 1104 37741
rect 869 37599 876 37655
rect 932 37599 1018 37655
rect 1074 37599 1104 37655
rect 869 37513 1104 37599
rect 3427 38142 3503 38154
rect 869 37457 876 37513
rect 932 37457 1018 37513
rect 1074 37457 1104 37513
rect 869 37371 1104 37457
rect 869 37315 876 37371
rect 932 37315 1018 37371
rect 1074 37315 1104 37371
rect 869 37229 1104 37315
rect 869 37173 876 37229
rect 932 37173 1018 37229
rect 1074 37173 1104 37229
rect 869 37154 1104 37173
rect 704 37087 1104 37154
rect 704 37031 734 37087
rect 790 37031 876 37087
rect 932 37031 1018 37087
rect 1074 37031 1104 37087
rect 704 36945 1104 37031
rect 704 36889 734 36945
rect 790 36889 876 36945
rect 932 36889 1018 36945
rect 1074 36889 1104 36945
rect 704 36803 1104 36889
rect 704 36747 734 36803
rect 790 36747 876 36803
rect 932 36747 1018 36803
rect 1074 36747 1104 36803
rect 704 36661 1104 36747
rect 704 36605 734 36661
rect 790 36605 876 36661
rect 932 36605 1018 36661
rect 1074 36605 1104 36661
rect 704 36519 1104 36605
rect 704 36463 734 36519
rect 790 36463 876 36519
rect 932 36463 1018 36519
rect 1074 36463 1104 36519
rect 704 36430 1104 36463
rect 2393 37569 2783 37581
rect 2393 37413 2719 37569
rect 2771 37413 2783 37569
rect 2393 37401 2783 37413
rect 3195 37569 3271 37581
rect 3195 37413 3207 37569
rect 3259 37413 3271 37569
rect 2393 36268 2469 37401
rect 2066 36256 2469 36268
rect 165 36178 383 36230
rect 165 36122 175 36178
rect 231 36122 317 36178
rect 373 36122 383 36178
rect 2066 36204 2088 36256
rect 2452 36204 2469 36256
rect 2066 36192 2469 36204
rect 165 36036 383 36122
rect 165 35980 175 36036
rect 231 35980 317 36036
rect 373 35980 383 36036
rect 165 35894 383 35980
rect 165 35838 175 35894
rect 231 35838 317 35894
rect 373 35838 383 35894
rect 1822 36120 2002 36132
rect 1822 36068 1834 36120
rect 1990 36068 2002 36120
rect 1822 36056 2002 36068
rect 165 35752 383 35838
rect 165 35696 175 35752
rect 231 35696 317 35752
rect 373 35696 383 35752
rect 165 35610 383 35696
rect 1310 35848 1490 35860
rect 1310 35796 1322 35848
rect 1478 35796 1490 35848
rect 1310 35784 1490 35796
rect 165 35554 175 35610
rect 231 35554 317 35610
rect 373 35554 383 35610
rect 165 35468 383 35554
rect 165 35412 175 35468
rect 231 35412 317 35468
rect 373 35412 383 35468
rect 165 35326 383 35412
rect 165 35270 175 35326
rect 231 35270 317 35326
rect 373 35270 383 35326
rect 165 35184 383 35270
rect 165 35128 175 35184
rect 231 35128 317 35184
rect 373 35128 383 35184
rect 165 35042 383 35128
rect 165 34986 175 35042
rect 231 34986 317 35042
rect 373 34986 383 35042
rect 165 34900 383 34986
rect 165 34844 175 34900
rect 231 34844 317 34900
rect 373 34844 383 34900
rect 165 34758 383 34844
rect 165 34702 175 34758
rect 231 34702 317 34758
rect 373 34702 383 34758
rect 165 34616 383 34702
rect 165 34560 175 34616
rect 231 34560 317 34616
rect 373 34560 383 34616
rect 165 34474 383 34560
rect 165 34418 175 34474
rect 231 34418 317 34474
rect 373 34418 383 34474
rect 165 34332 383 34418
rect 165 34276 175 34332
rect 231 34276 317 34332
rect 373 34276 383 34332
rect 165 34190 383 34276
rect 165 34134 175 34190
rect 231 34134 317 34190
rect 373 34134 383 34190
rect 165 34048 383 34134
rect 165 33992 175 34048
rect 231 33992 317 34048
rect 373 33992 383 34048
rect 165 33906 383 33992
rect 165 33850 175 33906
rect 231 33850 317 33906
rect 373 33850 383 33906
rect 165 33764 383 33850
rect 165 33708 175 33764
rect 231 33708 317 33764
rect 373 33708 383 33764
rect 165 33622 383 33708
rect 486 35617 562 35627
rect 486 35561 496 35617
rect 552 35561 562 35617
rect 486 35475 498 35561
rect 550 35475 562 35561
rect 486 35419 496 35475
rect 552 35419 562 35475
rect 486 35333 498 35419
rect 550 35333 562 35419
rect 486 35277 496 35333
rect 552 35277 562 35333
rect 486 35191 498 35277
rect 550 35191 562 35277
rect 486 35135 496 35191
rect 552 35135 562 35191
rect 486 35049 498 35135
rect 550 35049 562 35135
rect 486 34993 496 35049
rect 552 34993 562 35049
rect 486 34907 498 34993
rect 550 34907 562 34993
rect 486 34851 496 34907
rect 552 34851 562 34907
rect 486 34765 498 34851
rect 550 34765 562 34851
rect 486 34709 496 34765
rect 552 34709 562 34765
rect 486 34623 498 34709
rect 550 34623 562 34709
rect 486 34567 496 34623
rect 552 34567 562 34623
rect 486 34481 498 34567
rect 550 34481 562 34567
rect 486 34425 496 34481
rect 552 34425 562 34481
rect 486 34339 498 34425
rect 550 34339 562 34425
rect 486 34283 496 34339
rect 552 34283 562 34339
rect 486 34197 498 34283
rect 550 34197 562 34283
rect 486 34141 496 34197
rect 552 34141 562 34197
rect 486 34055 498 34141
rect 550 34055 562 34141
rect 724 35612 800 35622
rect 724 35556 734 35612
rect 790 35556 800 35612
rect 724 35470 736 35556
rect 788 35470 800 35556
rect 724 35414 734 35470
rect 790 35414 800 35470
rect 724 35328 736 35414
rect 788 35328 800 35414
rect 724 35272 734 35328
rect 790 35272 800 35328
rect 724 35186 736 35272
rect 788 35186 800 35272
rect 724 35130 734 35186
rect 790 35130 800 35186
rect 724 35044 736 35130
rect 788 35044 800 35130
rect 724 34988 734 35044
rect 790 34988 800 35044
rect 724 34902 736 34988
rect 788 34902 800 34988
rect 724 34846 734 34902
rect 790 34846 800 34902
rect 724 34760 736 34846
rect 788 34760 800 34846
rect 724 34704 734 34760
rect 790 34704 800 34760
rect 724 34618 736 34704
rect 788 34618 800 34704
rect 724 34562 734 34618
rect 790 34562 800 34618
rect 724 34476 736 34562
rect 788 34476 800 34562
rect 724 34420 734 34476
rect 790 34420 800 34476
rect 724 34334 736 34420
rect 788 34334 800 34420
rect 724 34278 734 34334
rect 790 34278 800 34334
rect 724 34192 736 34278
rect 788 34192 800 34278
rect 724 34136 734 34192
rect 790 34136 800 34192
rect 724 34126 800 34136
rect 486 33999 496 34055
rect 552 33999 562 34055
rect 486 33913 498 33999
rect 550 33913 562 33999
rect 486 33857 496 33913
rect 552 33857 562 33913
rect 486 33771 498 33857
rect 550 33771 562 33857
rect 486 33715 496 33771
rect 552 33715 562 33771
rect 486 33705 562 33715
rect 165 33566 175 33622
rect 231 33566 317 33622
rect 373 33566 383 33622
rect 165 33480 383 33566
rect 165 33424 175 33480
rect 231 33424 317 33480
rect 373 33424 383 33480
rect 165 33338 383 33424
rect 165 33282 175 33338
rect 231 33282 317 33338
rect 373 33282 383 33338
rect 165 28262 383 33282
rect 486 33481 562 33493
rect 486 32978 498 33481
rect 550 32978 562 33481
rect 486 32922 496 32978
rect 552 32922 562 32978
rect 486 32836 498 32922
rect 550 32836 562 32922
rect 486 32780 496 32836
rect 552 32780 562 32836
rect 486 32694 498 32780
rect 550 32694 562 32780
rect 486 32638 496 32694
rect 552 32638 562 32694
rect 486 32552 498 32638
rect 550 32552 562 32638
rect 486 32496 496 32552
rect 552 32496 562 32552
rect 1310 32518 1386 35784
rect 1822 34065 1898 36056
rect 1822 33909 1834 34065
rect 1886 33909 1898 34065
rect 1822 33897 1898 33909
rect 2066 34065 2142 36192
rect 3195 36132 3271 37413
rect 3091 36120 3271 36132
rect 3091 36068 3103 36120
rect 3259 36068 3271 36120
rect 3091 36056 3271 36068
rect 3427 37154 3439 38142
rect 3491 37154 3503 38142
rect 6049 38142 6125 38154
rect 6049 37797 6061 38142
rect 6113 37797 6125 38142
rect 6049 37741 6059 37797
rect 6115 37741 6125 37797
rect 6049 37655 6061 37741
rect 6113 37655 6125 37741
rect 6049 37599 6059 37655
rect 6115 37599 6125 37655
rect 2066 33909 2078 34065
rect 2130 33909 2142 34065
rect 2066 33897 2142 33909
rect 2482 35984 2662 35996
rect 2482 35932 2494 35984
rect 2650 35932 2662 35984
rect 2482 35920 2662 35932
rect 2482 34065 2558 35920
rect 3427 35860 3503 37154
rect 3659 37569 3735 37581
rect 3659 37413 3671 37569
rect 3723 37413 3735 37569
rect 3659 36132 3735 37413
rect 4147 37569 4537 37581
rect 4147 37413 4159 37569
rect 4211 37413 4537 37569
rect 4147 37401 4537 37413
rect 4461 36268 4537 37401
rect 6049 37513 6061 37599
rect 6113 37513 6125 37599
rect 6049 37457 6059 37513
rect 6115 37457 6125 37513
rect 6049 37371 6061 37457
rect 6113 37371 6125 37457
rect 6049 37315 6059 37371
rect 6115 37315 6125 37371
rect 6049 37229 6061 37315
rect 6113 37229 6125 37315
rect 6049 37173 6059 37229
rect 6115 37173 6125 37229
rect 6049 37154 6061 37173
rect 6113 37154 6125 37173
rect 6049 37087 6125 37154
rect 6049 37031 6059 37087
rect 6115 37031 6125 37087
rect 6049 36945 6125 37031
rect 6049 36889 6059 36945
rect 6115 36889 6125 36945
rect 6049 36803 6125 36889
rect 6049 36747 6059 36803
rect 6115 36747 6125 36803
rect 6049 36661 6125 36747
rect 6049 36605 6059 36661
rect 6115 36605 6125 36661
rect 6049 36519 6125 36605
rect 6049 36463 6059 36519
rect 6115 36463 6125 36519
rect 6049 36453 6125 36463
rect 4461 36256 4641 36268
rect 4461 36204 4473 36256
rect 4629 36204 4641 36256
rect 4461 36192 4641 36204
rect 5810 36256 5990 36268
rect 5810 36204 5822 36256
rect 5978 36204 5990 36256
rect 5810 36192 5990 36204
rect 3659 36120 3839 36132
rect 3659 36068 3671 36120
rect 3827 36068 3839 36120
rect 3659 36056 3839 36068
rect 5394 35984 5574 35996
rect 5394 35932 5406 35984
rect 5562 35932 5574 35984
rect 5394 35920 5574 35932
rect 3092 35784 3503 35860
rect 3092 35612 3168 35784
rect 3092 35556 3102 35612
rect 3158 35556 3168 35612
rect 3092 35470 3104 35556
rect 3156 35470 3168 35556
rect 3092 35414 3102 35470
rect 3158 35414 3168 35470
rect 3092 35328 3104 35414
rect 3156 35328 3168 35414
rect 3092 35272 3102 35328
rect 3158 35272 3168 35328
rect 3092 35186 3104 35272
rect 3156 35186 3168 35272
rect 3092 35130 3102 35186
rect 3158 35130 3168 35186
rect 3092 35044 3104 35130
rect 3156 35044 3168 35130
rect 3092 34988 3102 35044
rect 3158 34988 3168 35044
rect 3092 34902 3104 34988
rect 3156 34902 3168 34988
rect 3092 34846 3102 34902
rect 3158 34846 3168 34902
rect 3092 34760 3104 34846
rect 3156 34760 3168 34846
rect 3092 34704 3102 34760
rect 3158 34704 3168 34760
rect 3092 34618 3104 34704
rect 3156 34618 3168 34704
rect 3092 34562 3102 34618
rect 3158 34562 3168 34618
rect 3092 34476 3104 34562
rect 3156 34476 3168 34562
rect 3092 34420 3102 34476
rect 3158 34420 3168 34476
rect 3092 34334 3104 34420
rect 3156 34334 3168 34420
rect 3092 34278 3102 34334
rect 3158 34278 3168 34334
rect 3092 34192 3104 34278
rect 3156 34192 3168 34278
rect 3092 34136 3102 34192
rect 3158 34136 3168 34192
rect 3092 34126 3168 34136
rect 3386 35712 3566 35724
rect 3386 35660 3398 35712
rect 3554 35660 3566 35712
rect 3386 35648 3566 35660
rect 3990 35716 4066 35726
rect 3990 35660 4000 35716
rect 4056 35660 4066 35716
rect 2482 33909 2494 34065
rect 2546 33909 2558 34065
rect 2482 33897 2558 33909
rect 3386 33897 3462 35648
rect 3990 35576 4066 35660
rect 4490 35712 4670 35724
rect 4490 35660 4502 35712
rect 4658 35660 4670 35712
rect 4490 35648 4670 35660
rect 3990 35574 4002 35576
rect 4054 35574 4066 35576
rect 3990 35518 4000 35574
rect 4056 35518 4066 35574
rect 3990 35432 4002 35518
rect 4054 35432 4066 35518
rect 3990 35376 4000 35432
rect 4056 35376 4066 35432
rect 3990 35290 4002 35376
rect 4054 35290 4066 35376
rect 3990 35234 4000 35290
rect 4056 35234 4066 35290
rect 3990 35148 4002 35234
rect 4054 35148 4066 35234
rect 3990 35092 4000 35148
rect 4056 35092 4066 35148
rect 3990 35006 4002 35092
rect 4054 35006 4066 35092
rect 3990 34950 4000 35006
rect 4056 34950 4066 35006
rect 3990 34864 4002 34950
rect 4054 34864 4066 34950
rect 3990 34808 4000 34864
rect 4056 34808 4066 34864
rect 3990 34722 4002 34808
rect 4054 34722 4066 34808
rect 3990 34666 4000 34722
rect 4056 34666 4066 34722
rect 3990 34580 4002 34666
rect 4054 34580 4066 34666
rect 3990 34524 4000 34580
rect 4056 34524 4066 34580
rect 3990 34438 4002 34524
rect 4054 34438 4066 34524
rect 3990 34382 4000 34438
rect 4056 34382 4066 34438
rect 3990 34296 4002 34382
rect 4054 34296 4066 34382
rect 3990 34240 4000 34296
rect 4056 34240 4066 34296
rect 3990 34154 4002 34240
rect 4054 34154 4066 34240
rect 3990 34098 4000 34154
rect 4056 34098 4066 34154
rect 3990 34012 4002 34098
rect 4054 34012 4066 34098
rect 3990 33956 4000 34012
rect 4056 33956 4066 34012
rect 3990 33870 4002 33956
rect 4054 33870 4066 33956
rect 4594 33897 4670 35648
rect 4888 35612 4964 35622
rect 4888 35556 4898 35612
rect 4954 35556 4964 35612
rect 4888 35470 4900 35556
rect 4952 35470 4964 35556
rect 4888 35414 4898 35470
rect 4954 35414 4964 35470
rect 4888 35328 4900 35414
rect 4952 35328 4964 35414
rect 4888 35272 4898 35328
rect 4954 35272 4964 35328
rect 4888 35186 4900 35272
rect 4952 35186 4964 35272
rect 4888 35130 4898 35186
rect 4954 35130 4964 35186
rect 4888 35044 4900 35130
rect 4952 35044 4964 35130
rect 4888 34988 4898 35044
rect 4954 34988 4964 35044
rect 4888 34902 4900 34988
rect 4952 34902 4964 34988
rect 4888 34846 4898 34902
rect 4954 34846 4964 34902
rect 4888 34760 4900 34846
rect 4952 34760 4964 34846
rect 4888 34704 4898 34760
rect 4954 34704 4964 34760
rect 4888 34618 4900 34704
rect 4952 34618 4964 34704
rect 4888 34562 4898 34618
rect 4954 34562 4964 34618
rect 4888 34476 4900 34562
rect 4952 34476 4964 34562
rect 4888 34420 4898 34476
rect 4954 34420 4964 34476
rect 4888 34334 4900 34420
rect 4952 34334 4964 34420
rect 4888 34278 4898 34334
rect 4954 34278 4964 34334
rect 4888 34192 4900 34278
rect 4952 34192 4964 34278
rect 4888 34136 4898 34192
rect 4954 34136 4964 34192
rect 4888 34126 4964 34136
rect 5498 34065 5574 35920
rect 5498 33909 5510 34065
rect 5562 33909 5574 34065
rect 5498 33897 5574 33909
rect 5914 34065 5990 36192
rect 6054 36120 6234 36132
rect 6054 36068 6066 36120
rect 6222 36068 6234 36120
rect 6054 36056 6234 36068
rect 5914 33909 5926 34065
rect 5978 33909 5990 34065
rect 5914 33897 5990 33909
rect 6158 34065 6234 36056
rect 6566 35848 6746 35860
rect 6566 35796 6578 35848
rect 6734 35796 6746 35848
rect 6566 35784 6746 35796
rect 6158 33909 6170 34065
rect 6222 33909 6234 34065
rect 6158 33897 6234 33909
rect 3990 33814 4000 33870
rect 4056 33814 4066 33870
rect 3990 33728 4002 33814
rect 4054 33728 4066 33814
rect 3990 33672 4000 33728
rect 4056 33672 4066 33728
rect 3990 33586 4002 33672
rect 4054 33586 4066 33672
rect 3990 33530 4000 33586
rect 4056 33530 4066 33586
rect 3990 33444 4002 33530
rect 4054 33444 4066 33530
rect 3990 33388 4000 33444
rect 4056 33388 4066 33444
rect 3990 33302 4002 33388
rect 4054 33302 4066 33388
rect 3990 33246 4000 33302
rect 4056 33246 4066 33302
rect 3990 32924 4002 33246
rect 4054 32924 4066 33246
rect 3990 32912 4066 32924
rect 3990 32535 4066 32545
rect 486 32410 498 32496
rect 550 32410 562 32496
rect 486 32354 496 32410
rect 552 32354 562 32410
rect 486 32268 498 32354
rect 550 32268 562 32354
rect 3990 32479 4000 32535
rect 4056 32479 4066 32535
rect 6670 32518 6746 35784
rect 3990 32455 4066 32479
rect 3990 32393 4002 32455
rect 4054 32393 4066 32455
rect 3990 32337 4000 32393
rect 4056 32337 4066 32393
rect 486 32212 496 32268
rect 552 32212 562 32268
rect 486 32126 498 32212
rect 550 32126 562 32212
rect 486 32070 496 32126
rect 552 32070 562 32126
rect 486 31984 498 32070
rect 550 31984 562 32070
rect 486 31928 496 31984
rect 552 31928 562 31984
rect 486 31842 498 31928
rect 550 31842 562 31928
rect 486 31786 496 31842
rect 552 31786 562 31842
rect 486 31700 498 31786
rect 550 31700 562 31786
rect 486 31644 496 31700
rect 552 31644 562 31700
rect 486 31558 498 31644
rect 550 31558 562 31644
rect 486 31502 496 31558
rect 552 31502 562 31558
rect 486 31416 498 31502
rect 550 31416 562 31502
rect 486 31360 496 31416
rect 552 31360 562 31416
rect 486 31274 498 31360
rect 550 31274 562 31360
rect 486 31218 496 31274
rect 552 31218 562 31274
rect 486 31132 498 31218
rect 550 31132 562 31218
rect 486 31076 496 31132
rect 552 31076 562 31132
rect 486 30990 498 31076
rect 550 30990 562 31076
rect 486 30934 496 30990
rect 552 30934 562 30990
rect 486 30848 498 30934
rect 550 30848 562 30934
rect 486 30792 496 30848
rect 552 30792 562 30848
rect 486 30706 498 30792
rect 550 30706 562 30792
rect 486 30650 496 30706
rect 552 30650 562 30706
rect 486 30564 498 30650
rect 550 30564 562 30650
rect 486 30508 496 30564
rect 552 30508 562 30564
rect 486 30422 498 30508
rect 550 30422 562 30508
rect 486 30366 496 30422
rect 552 30366 562 30422
rect 486 30280 498 30366
rect 550 30280 562 30366
rect 486 30224 496 30280
rect 552 30224 562 30280
rect 486 30138 498 30224
rect 550 30138 562 30224
rect 486 30082 496 30138
rect 552 30082 562 30138
rect 486 29685 498 30082
rect 550 29685 562 30082
rect 968 32322 1044 32332
rect 968 32266 978 32322
rect 1034 32266 1044 32322
rect 968 32180 980 32266
rect 1032 32180 1044 32266
rect 968 32124 978 32180
rect 1034 32124 1044 32180
rect 968 32038 980 32124
rect 1032 32038 1044 32124
rect 968 31982 978 32038
rect 1034 31982 1044 32038
rect 968 31896 980 31982
rect 1032 31896 1044 31982
rect 968 31840 978 31896
rect 1034 31840 1044 31896
rect 968 31754 980 31840
rect 1032 31754 1044 31840
rect 968 31698 978 31754
rect 1034 31698 1044 31754
rect 968 31612 980 31698
rect 1032 31612 1044 31698
rect 968 31556 978 31612
rect 1034 31556 1044 31612
rect 968 31470 980 31556
rect 1032 31470 1044 31556
rect 968 31414 978 31470
rect 1034 31414 1044 31470
rect 968 31328 980 31414
rect 1032 31328 1044 31414
rect 968 31272 978 31328
rect 1034 31272 1044 31328
rect 968 31186 980 31272
rect 1032 31186 1044 31272
rect 968 31130 978 31186
rect 1034 31130 1044 31186
rect 968 31044 980 31130
rect 1032 31044 1044 31130
rect 968 30988 978 31044
rect 1034 30988 1044 31044
rect 968 30902 980 30988
rect 1032 30902 1044 30988
rect 968 30846 978 30902
rect 1034 30846 1044 30902
rect 968 30760 980 30846
rect 1032 30760 1044 30846
rect 968 30704 978 30760
rect 1034 30704 1044 30760
rect 968 30618 980 30704
rect 1032 30618 1044 30704
rect 968 30562 978 30618
rect 1034 30562 1044 30618
rect 968 30476 980 30562
rect 1032 30476 1044 30562
rect 968 30420 978 30476
rect 1034 30420 1044 30476
rect 968 30334 980 30420
rect 1032 30334 1044 30420
rect 968 30278 978 30334
rect 1034 30278 1044 30334
rect 2360 32322 2436 32332
rect 2360 32266 2370 32322
rect 2426 32266 2436 32322
rect 2360 32180 2372 32266
rect 2424 32180 2436 32266
rect 2360 32124 2370 32180
rect 2426 32124 2436 32180
rect 2360 32038 2372 32124
rect 2424 32038 2436 32124
rect 2360 31982 2370 32038
rect 2426 31982 2436 32038
rect 2360 31896 2372 31982
rect 2424 31896 2436 31982
rect 2360 31840 2370 31896
rect 2426 31840 2436 31896
rect 2360 31754 2372 31840
rect 2424 31754 2436 31840
rect 2360 31698 2370 31754
rect 2426 31698 2436 31754
rect 2360 31612 2372 31698
rect 2424 31612 2436 31698
rect 2360 31556 2370 31612
rect 2426 31556 2436 31612
rect 2360 31470 2372 31556
rect 2424 31470 2436 31556
rect 2360 31414 2370 31470
rect 2426 31414 2436 31470
rect 2360 31328 2372 31414
rect 2424 31328 2436 31414
rect 2360 31272 2370 31328
rect 2426 31272 2436 31328
rect 2360 31186 2372 31272
rect 2424 31186 2436 31272
rect 2360 31130 2370 31186
rect 2426 31130 2436 31186
rect 2360 31044 2372 31130
rect 2424 31044 2436 31130
rect 2360 30988 2370 31044
rect 2426 30988 2436 31044
rect 2360 30902 2372 30988
rect 2424 30902 2436 30988
rect 2360 30846 2370 30902
rect 2426 30846 2436 30902
rect 2360 30760 2372 30846
rect 2424 30760 2436 30846
rect 2360 30704 2370 30760
rect 2426 30704 2436 30760
rect 2360 30618 2372 30704
rect 2424 30618 2436 30704
rect 2360 30562 2370 30618
rect 2426 30562 2436 30618
rect 2360 30476 2372 30562
rect 2424 30476 2436 30562
rect 2360 30420 2370 30476
rect 2426 30420 2436 30476
rect 2360 30334 2372 30420
rect 2424 30334 2436 30420
rect 968 30192 980 30278
rect 1032 30192 1044 30278
rect 968 30136 978 30192
rect 1034 30136 1044 30192
rect 968 30084 980 30136
rect 1032 30084 1044 30136
rect 968 30072 1044 30084
rect 1444 30308 1544 30320
rect 1444 29944 1468 30308
rect 1520 29944 1544 30308
rect 1444 29831 1544 29944
rect 486 29673 562 29685
rect 1007 29731 1544 29831
rect 1688 30308 1788 30320
rect 1688 29944 1712 30308
rect 1764 29944 1788 30308
rect 2360 30278 2370 30334
rect 2426 30278 2436 30334
rect 2360 30192 2372 30278
rect 2424 30192 2436 30278
rect 2360 30136 2370 30192
rect 2426 30136 2436 30192
rect 2360 30084 2372 30136
rect 2424 30084 2436 30136
rect 2360 30072 2436 30084
rect 2776 32322 2852 32332
rect 2776 32266 2786 32322
rect 2842 32266 2852 32322
rect 2776 32180 2788 32266
rect 2840 32180 2852 32266
rect 2776 32124 2786 32180
rect 2842 32124 2852 32180
rect 2776 32038 2788 32124
rect 2840 32038 2852 32124
rect 2776 31982 2786 32038
rect 2842 31982 2852 32038
rect 2776 31896 2788 31982
rect 2840 31896 2852 31982
rect 2776 31840 2786 31896
rect 2842 31840 2852 31896
rect 2776 31754 2788 31840
rect 2840 31754 2852 31840
rect 2776 31698 2786 31754
rect 2842 31698 2852 31754
rect 2776 31612 2788 31698
rect 2840 31612 2852 31698
rect 2776 31556 2786 31612
rect 2842 31556 2852 31612
rect 2776 31470 2788 31556
rect 2840 31470 2852 31556
rect 2776 31414 2786 31470
rect 2842 31414 2852 31470
rect 2776 31328 2788 31414
rect 2840 31328 2852 31414
rect 2776 31272 2786 31328
rect 2842 31272 2852 31328
rect 2776 31186 2788 31272
rect 2840 31186 2852 31272
rect 2776 31130 2786 31186
rect 2842 31130 2852 31186
rect 2776 31044 2788 31130
rect 2840 31044 2852 31130
rect 2776 30988 2786 31044
rect 2842 30988 2852 31044
rect 2776 30902 2788 30988
rect 2840 30902 2852 30988
rect 2776 30846 2786 30902
rect 2842 30846 2852 30902
rect 2776 30760 2788 30846
rect 2840 30760 2852 30846
rect 2776 30704 2786 30760
rect 2842 30704 2852 30760
rect 2776 30618 2788 30704
rect 2840 30618 2852 30704
rect 3264 32323 3340 32333
rect 3264 32267 3274 32323
rect 3330 32267 3340 32323
rect 3264 32181 3276 32267
rect 3328 32181 3340 32267
rect 3264 32125 3274 32181
rect 3330 32125 3340 32181
rect 3264 32039 3276 32125
rect 3328 32039 3340 32125
rect 3264 31983 3274 32039
rect 3330 31983 3340 32039
rect 3264 31897 3276 31983
rect 3328 31897 3340 31983
rect 3264 31841 3274 31897
rect 3330 31841 3340 31897
rect 3264 31755 3276 31841
rect 3328 31755 3340 31841
rect 3264 31699 3274 31755
rect 3330 31699 3340 31755
rect 3264 31613 3276 31699
rect 3328 31613 3340 31699
rect 3264 31557 3274 31613
rect 3330 31557 3340 31613
rect 3264 31471 3276 31557
rect 3328 31471 3340 31557
rect 3264 31415 3274 31471
rect 3330 31415 3340 31471
rect 3264 31329 3276 31415
rect 3328 31329 3340 31415
rect 3264 31273 3274 31329
rect 3330 31273 3340 31329
rect 3264 31187 3276 31273
rect 3328 31187 3340 31273
rect 3264 31131 3274 31187
rect 3330 31131 3340 31187
rect 3264 31045 3276 31131
rect 3328 31045 3340 31131
rect 3264 30989 3274 31045
rect 3330 30989 3340 31045
rect 3264 30903 3276 30989
rect 3328 30903 3340 30989
rect 3264 30847 3274 30903
rect 3330 30847 3340 30903
rect 3264 30761 3276 30847
rect 3328 30761 3340 30847
rect 3264 30705 3274 30761
rect 3330 30705 3340 30761
rect 3264 30695 3340 30705
rect 3752 32272 3828 32282
rect 3752 32216 3762 32272
rect 3818 32216 3828 32272
rect 3752 32130 3764 32216
rect 3816 32130 3828 32216
rect 3752 32074 3762 32130
rect 3818 32074 3828 32130
rect 3752 31988 3764 32074
rect 3816 31988 3828 32074
rect 3752 31932 3762 31988
rect 3818 31932 3828 31988
rect 3752 31846 3764 31932
rect 3816 31846 3828 31932
rect 3752 31790 3762 31846
rect 3818 31790 3828 31846
rect 3752 31704 3764 31790
rect 3816 31704 3828 31790
rect 3752 31648 3762 31704
rect 3818 31648 3828 31704
rect 3752 31562 3764 31648
rect 3816 31562 3828 31648
rect 3752 31506 3762 31562
rect 3818 31506 3828 31562
rect 3752 31420 3764 31506
rect 3816 31420 3828 31506
rect 3752 31364 3762 31420
rect 3818 31364 3828 31420
rect 3752 31278 3764 31364
rect 3816 31278 3828 31364
rect 3752 31222 3762 31278
rect 3818 31222 3828 31278
rect 3752 31136 3764 31222
rect 3816 31136 3828 31222
rect 3752 31080 3762 31136
rect 3818 31080 3828 31136
rect 3752 30994 3764 31080
rect 3816 30994 3828 31080
rect 3752 30938 3762 30994
rect 3818 30938 3828 30994
rect 3752 30852 3764 30938
rect 3816 30852 3828 30938
rect 3752 30796 3762 30852
rect 3818 30796 3828 30852
rect 3752 30710 3764 30796
rect 3816 30710 3828 30796
rect 3752 30654 3762 30710
rect 3818 30654 3828 30710
rect 3752 30644 3828 30654
rect 3990 32251 4002 32337
rect 4054 32251 4066 32337
rect 4716 32323 4792 32333
rect 3990 32195 4000 32251
rect 4056 32195 4066 32251
rect 3990 32109 4002 32195
rect 4054 32109 4066 32195
rect 3990 32053 4000 32109
rect 4056 32053 4066 32109
rect 3990 31967 4002 32053
rect 4054 31967 4066 32053
rect 3990 31911 4000 31967
rect 4056 31911 4066 31967
rect 3990 31825 4002 31911
rect 4054 31825 4066 31911
rect 3990 31769 4000 31825
rect 4056 31769 4066 31825
rect 3990 31683 4002 31769
rect 4054 31683 4066 31769
rect 3990 31627 4000 31683
rect 4056 31627 4066 31683
rect 3990 31541 4002 31627
rect 4054 31541 4066 31627
rect 3990 31485 4000 31541
rect 4056 31485 4066 31541
rect 3990 31399 4002 31485
rect 4054 31399 4066 31485
rect 3990 31343 4000 31399
rect 4056 31343 4066 31399
rect 3990 31257 4002 31343
rect 4054 31257 4066 31343
rect 3990 31201 4000 31257
rect 4056 31201 4066 31257
rect 3990 31115 4002 31201
rect 4054 31115 4066 31201
rect 3990 31059 4000 31115
rect 4056 31059 4066 31115
rect 3990 30973 4002 31059
rect 4054 30973 4066 31059
rect 3990 30917 4000 30973
rect 4056 30917 4066 30973
rect 3990 30831 4002 30917
rect 4054 30831 4066 30917
rect 3990 30775 4000 30831
rect 4056 30775 4066 30831
rect 3990 30689 4002 30775
rect 4054 30689 4066 30775
rect 3990 30633 4000 30689
rect 4056 30633 4066 30689
rect 4228 32272 4304 32282
rect 4228 32216 4238 32272
rect 4294 32216 4304 32272
rect 4228 32130 4240 32216
rect 4292 32130 4304 32216
rect 4228 32074 4238 32130
rect 4294 32074 4304 32130
rect 4228 31988 4240 32074
rect 4292 31988 4304 32074
rect 4228 31932 4238 31988
rect 4294 31932 4304 31988
rect 4228 31846 4240 31932
rect 4292 31846 4304 31932
rect 4228 31790 4238 31846
rect 4294 31790 4304 31846
rect 4228 31704 4240 31790
rect 4292 31704 4304 31790
rect 4228 31648 4238 31704
rect 4294 31648 4304 31704
rect 4228 31562 4240 31648
rect 4292 31562 4304 31648
rect 4228 31506 4238 31562
rect 4294 31506 4304 31562
rect 4228 31420 4240 31506
rect 4292 31420 4304 31506
rect 4228 31364 4238 31420
rect 4294 31364 4304 31420
rect 4228 31278 4240 31364
rect 4292 31278 4304 31364
rect 4228 31222 4238 31278
rect 4294 31222 4304 31278
rect 4228 31136 4240 31222
rect 4292 31136 4304 31222
rect 4228 31080 4238 31136
rect 4294 31080 4304 31136
rect 4228 30994 4240 31080
rect 4292 30994 4304 31080
rect 4228 30938 4238 30994
rect 4294 30938 4304 30994
rect 4228 30852 4240 30938
rect 4292 30852 4304 30938
rect 4228 30796 4238 30852
rect 4294 30796 4304 30852
rect 4228 30710 4240 30796
rect 4292 30710 4304 30796
rect 4228 30654 4238 30710
rect 4294 30654 4304 30710
rect 4716 32267 4726 32323
rect 4782 32267 4792 32323
rect 4716 32181 4728 32267
rect 4780 32181 4792 32267
rect 4716 32125 4726 32181
rect 4782 32125 4792 32181
rect 4716 32039 4728 32125
rect 4780 32039 4792 32125
rect 4716 31983 4726 32039
rect 4782 31983 4792 32039
rect 4716 31897 4728 31983
rect 4780 31897 4792 31983
rect 4716 31841 4726 31897
rect 4782 31841 4792 31897
rect 4716 31755 4728 31841
rect 4780 31755 4792 31841
rect 4716 31699 4726 31755
rect 4782 31699 4792 31755
rect 4716 31613 4728 31699
rect 4780 31613 4792 31699
rect 4716 31557 4726 31613
rect 4782 31557 4792 31613
rect 4716 31471 4728 31557
rect 4780 31471 4792 31557
rect 4716 31415 4726 31471
rect 4782 31415 4792 31471
rect 4716 31329 4728 31415
rect 4780 31329 4792 31415
rect 4716 31273 4726 31329
rect 4782 31273 4792 31329
rect 4716 31187 4728 31273
rect 4780 31187 4792 31273
rect 4716 31131 4726 31187
rect 4782 31131 4792 31187
rect 4716 31045 4728 31131
rect 4780 31045 4792 31131
rect 4716 30989 4726 31045
rect 4782 30989 4792 31045
rect 4716 30903 4728 30989
rect 4780 30903 4792 30989
rect 4716 30847 4726 30903
rect 4782 30847 4792 30903
rect 4716 30761 4728 30847
rect 4780 30761 4792 30847
rect 4716 30705 4726 30761
rect 4782 30705 4792 30761
rect 4716 30695 4792 30705
rect 5204 32323 5280 32333
rect 5204 32267 5214 32323
rect 5270 32267 5280 32323
rect 5204 32181 5216 32267
rect 5268 32181 5280 32267
rect 5204 32125 5214 32181
rect 5270 32125 5280 32181
rect 5204 32039 5216 32125
rect 5268 32039 5280 32125
rect 5204 31983 5214 32039
rect 5270 31983 5280 32039
rect 5204 31897 5216 31983
rect 5268 31897 5280 31983
rect 5204 31841 5214 31897
rect 5270 31841 5280 31897
rect 5204 31755 5216 31841
rect 5268 31755 5280 31841
rect 5204 31699 5214 31755
rect 5270 31699 5280 31755
rect 5204 31613 5216 31699
rect 5268 31613 5280 31699
rect 5204 31557 5214 31613
rect 5270 31557 5280 31613
rect 5204 31471 5216 31557
rect 5268 31471 5280 31557
rect 5204 31415 5214 31471
rect 5270 31415 5280 31471
rect 5204 31329 5216 31415
rect 5268 31329 5280 31415
rect 5204 31273 5214 31329
rect 5270 31273 5280 31329
rect 5204 31187 5216 31273
rect 5268 31187 5280 31273
rect 5204 31131 5214 31187
rect 5270 31131 5280 31187
rect 5204 31045 5216 31131
rect 5268 31045 5280 31131
rect 5204 30989 5214 31045
rect 5270 30989 5280 31045
rect 5204 30903 5216 30989
rect 5268 30903 5280 30989
rect 5204 30847 5214 30903
rect 5270 30847 5280 30903
rect 5204 30761 5216 30847
rect 5268 30761 5280 30847
rect 5204 30705 5214 30761
rect 5270 30705 5280 30761
rect 5204 30695 5280 30705
rect 5620 32323 5696 32333
rect 5620 32267 5630 32323
rect 5686 32267 5696 32323
rect 5620 32181 5632 32267
rect 5684 32181 5696 32267
rect 5620 32125 5630 32181
rect 5686 32125 5696 32181
rect 5620 32039 5632 32125
rect 5684 32039 5696 32125
rect 5620 31983 5630 32039
rect 5686 31983 5696 32039
rect 5620 31897 5632 31983
rect 5684 31897 5696 31983
rect 5620 31841 5630 31897
rect 5686 31841 5696 31897
rect 5620 31755 5632 31841
rect 5684 31755 5696 31841
rect 5620 31699 5630 31755
rect 5686 31699 5696 31755
rect 5620 31613 5632 31699
rect 5684 31613 5696 31699
rect 5620 31557 5630 31613
rect 5686 31557 5696 31613
rect 5620 31471 5632 31557
rect 5684 31471 5696 31557
rect 5620 31415 5630 31471
rect 5686 31415 5696 31471
rect 5620 31329 5632 31415
rect 5684 31329 5696 31415
rect 5620 31273 5630 31329
rect 5686 31273 5696 31329
rect 5620 31187 5632 31273
rect 5684 31187 5696 31273
rect 5620 31131 5630 31187
rect 5686 31131 5696 31187
rect 5620 31045 5632 31131
rect 5684 31045 5696 31131
rect 5620 30989 5630 31045
rect 5686 30989 5696 31045
rect 5620 30903 5632 30989
rect 5684 30903 5696 30989
rect 5620 30847 5630 30903
rect 5686 30847 5696 30903
rect 5620 30761 5632 30847
rect 5684 30761 5696 30847
rect 5620 30705 5630 30761
rect 5686 30705 5696 30761
rect 5620 30695 5696 30705
rect 7012 32322 7088 32332
rect 7012 32266 7022 32322
rect 7078 32266 7088 32322
rect 7012 32180 7024 32266
rect 7076 32180 7088 32266
rect 7012 32124 7022 32180
rect 7078 32124 7088 32180
rect 7012 32038 7024 32124
rect 7076 32038 7088 32124
rect 7012 31982 7022 32038
rect 7078 31982 7088 32038
rect 7012 31896 7024 31982
rect 7076 31896 7088 31982
rect 7012 31840 7022 31896
rect 7078 31840 7088 31896
rect 7012 31754 7024 31840
rect 7076 31754 7088 31840
rect 7012 31698 7022 31754
rect 7078 31698 7088 31754
rect 7012 31612 7024 31698
rect 7076 31612 7088 31698
rect 7012 31556 7022 31612
rect 7078 31556 7088 31612
rect 7012 31470 7024 31556
rect 7076 31470 7088 31556
rect 7012 31414 7022 31470
rect 7078 31414 7088 31470
rect 7012 31328 7024 31414
rect 7076 31328 7088 31414
rect 7012 31272 7022 31328
rect 7078 31272 7088 31328
rect 7012 31186 7024 31272
rect 7076 31186 7088 31272
rect 7012 31130 7022 31186
rect 7078 31130 7088 31186
rect 7012 31044 7024 31130
rect 7076 31044 7088 31130
rect 7012 30988 7022 31044
rect 7078 30988 7088 31044
rect 7012 30902 7024 30988
rect 7076 30902 7088 30988
rect 7012 30846 7022 30902
rect 7078 30846 7088 30902
rect 7012 30760 7024 30846
rect 7076 30760 7088 30846
rect 7012 30704 7022 30760
rect 7078 30704 7088 30760
rect 4228 30644 4304 30654
rect 3990 30623 4066 30633
rect 2776 30562 2786 30618
rect 2842 30562 2852 30618
rect 2776 30476 2788 30562
rect 2840 30476 2852 30562
rect 7012 30618 7024 30704
rect 7076 30618 7088 30704
rect 7012 30562 7022 30618
rect 7078 30562 7088 30618
rect 2776 30420 2786 30476
rect 2842 30420 2852 30476
rect 2776 30334 2788 30420
rect 2840 30334 2852 30420
rect 2776 30278 2786 30334
rect 2842 30278 2852 30334
rect 2776 30192 2788 30278
rect 2840 30192 2852 30278
rect 2776 30136 2786 30192
rect 2842 30136 2852 30192
rect 2776 30084 2788 30136
rect 2840 30084 2852 30136
rect 3020 30488 4243 30500
rect 3020 30124 3032 30488
rect 3084 30400 4243 30488
rect 3084 30124 3096 30400
rect 3020 30112 3096 30124
rect 3496 30308 3596 30320
rect 2776 30072 2852 30084
rect 165 28197 586 28262
rect 165 28141 175 28197
rect 231 28141 317 28197
rect 373 28141 586 28197
rect 165 28055 586 28141
rect 165 27999 175 28055
rect 231 27999 317 28055
rect 373 28005 586 28055
rect 1007 28031 1107 29731
rect 1688 29651 1788 29944
rect 3496 29944 3520 30308
rect 3572 29944 3596 30308
rect 1985 29739 3339 29749
rect 1985 29683 1995 29739
rect 2051 29737 2137 29739
rect 2193 29737 2279 29739
rect 2335 29737 2421 29739
rect 2477 29737 2563 29739
rect 2619 29737 2705 29739
rect 2761 29737 2847 29739
rect 2903 29737 2989 29739
rect 3045 29737 3131 29739
rect 3187 29737 3273 29739
rect 2051 29683 2137 29685
rect 2193 29683 2279 29685
rect 2335 29683 2421 29685
rect 2477 29683 2563 29685
rect 2619 29683 2705 29685
rect 2761 29683 2847 29685
rect 2903 29683 2989 29685
rect 3045 29683 3131 29685
rect 3187 29683 3273 29685
rect 3329 29683 3339 29739
rect 1985 29673 3339 29683
rect 1187 29551 1788 29651
rect 1187 28031 1287 29551
rect 1367 29447 1547 29459
rect 1367 29395 1379 29447
rect 1535 29395 1547 29447
rect 1367 29383 1547 29395
rect 1367 28031 1467 29383
rect 1547 29267 1727 29279
rect 1547 29215 1559 29267
rect 1715 29215 1727 29267
rect 1547 29203 1727 29215
rect 1547 28031 1655 29203
rect 3496 29072 3596 29944
rect 4143 29099 4243 30400
rect 4472 30488 6002 30500
rect 4472 30124 4484 30488
rect 4536 30400 6002 30488
rect 4536 30124 4548 30400
rect 4472 30112 4548 30124
rect 4948 30308 5048 30320
rect 3496 29060 3676 29072
rect 3496 29008 3508 29060
rect 3664 29008 3676 29060
rect 3496 28996 3676 29008
rect 4143 28943 4167 29099
rect 4219 28943 4243 29099
rect 4143 28931 4243 28943
rect 4948 29944 4972 30308
rect 5024 29944 5048 30308
rect 4948 29099 5048 29944
rect 4948 28943 4972 29099
rect 5024 28943 5048 29099
rect 4948 28931 5048 28943
rect 5902 29099 6002 30400
rect 7012 30476 7024 30562
rect 7076 30476 7088 30562
rect 7012 30420 7022 30476
rect 7078 30420 7088 30476
rect 7012 30334 7024 30420
rect 7076 30334 7088 30420
rect 6512 30308 6612 30320
rect 6512 29944 6536 30308
rect 6588 29944 6612 30308
rect 6512 29459 6612 29944
rect 6432 29447 6612 29459
rect 6432 29395 6444 29447
rect 6600 29395 6612 29447
rect 6432 29383 6612 29395
rect 6756 30308 6856 30320
rect 6756 29944 6780 30308
rect 6832 29944 6856 30308
rect 7012 30278 7022 30334
rect 7078 30278 7088 30334
rect 7012 30192 7024 30278
rect 7076 30192 7088 30278
rect 7012 30136 7022 30192
rect 7078 30136 7088 30192
rect 7012 30084 7024 30136
rect 7076 30084 7088 30136
rect 7012 30072 7088 30084
rect 6756 29279 6856 29944
rect 6676 29267 6856 29279
rect 6676 29215 6688 29267
rect 6844 29215 6856 29267
rect 6676 29203 6856 29215
rect 5902 28943 5926 29099
rect 5978 28943 6002 29099
rect 5902 28931 6002 28943
rect 373 27999 383 28005
rect 165 27913 383 27999
rect 165 27857 175 27913
rect 231 27857 317 27913
rect 373 27857 383 27913
rect 165 27771 383 27857
rect 165 27715 175 27771
rect 231 27715 317 27771
rect 373 27715 383 27771
rect 165 27629 383 27715
rect 7332 27675 7732 41308
rect 11356 41288 11517 41444
rect 11569 41288 11581 41444
rect 11356 41276 11581 41288
rect 11137 40793 11213 40805
rect 11137 40637 11149 40793
rect 11201 40637 11213 40793
rect 11356 40730 11432 41276
rect 11520 40971 12060 40983
rect 11520 40815 11532 40971
rect 11584 40815 12060 40971
rect 11520 40803 12060 40815
rect 11356 40654 11596 40730
rect 11137 40514 11213 40637
rect 11137 40438 11276 40514
rect 10784 40364 10964 40376
rect 10784 40312 10796 40364
rect 10952 40312 10964 40364
rect 10784 40300 10964 40312
rect 10644 40092 10824 40104
rect 10644 40040 10656 40092
rect 10812 40040 10824 40092
rect 10644 40028 10824 40040
rect 7888 39946 9767 39956
rect 7888 39944 7997 39946
rect 8053 39944 8139 39946
rect 8195 39944 8281 39946
rect 8337 39944 8423 39946
rect 8479 39944 8565 39946
rect 8621 39944 8707 39946
rect 8763 39944 8849 39946
rect 8905 39944 8991 39946
rect 9047 39944 9133 39946
rect 9189 39944 9275 39946
rect 9331 39944 9417 39946
rect 9473 39944 9559 39946
rect 9615 39944 9701 39946
rect 7888 39892 7900 39944
rect 7888 39890 7997 39892
rect 8053 39890 8139 39892
rect 8195 39890 8281 39892
rect 8337 39890 8423 39892
rect 8479 39890 8565 39892
rect 8621 39890 8707 39892
rect 8763 39890 8849 39892
rect 8905 39890 8991 39892
rect 9047 39890 9133 39892
rect 9189 39890 9275 39892
rect 9331 39890 9417 39892
rect 9473 39890 9559 39892
rect 9615 39890 9701 39892
rect 9757 39890 9767 39946
rect 7888 39880 9767 39890
rect 10327 39418 10403 39430
rect 10327 39414 10339 39418
rect 10391 39414 10403 39418
rect 10327 39358 10337 39414
rect 10393 39358 10403 39414
rect 10327 39272 10339 39358
rect 10391 39272 10403 39358
rect 10327 39216 10337 39272
rect 10393 39216 10403 39272
rect 10327 39130 10339 39216
rect 10391 39130 10403 39216
rect 10327 39074 10337 39130
rect 10393 39074 10403 39130
rect 10327 38988 10339 39074
rect 10391 38988 10403 39074
rect 10327 38932 10337 38988
rect 10393 38932 10403 38988
rect 10327 38846 10339 38932
rect 10391 38846 10403 38932
rect 10327 38790 10337 38846
rect 10393 38790 10403 38846
rect 10327 38704 10339 38790
rect 10391 38704 10403 38790
rect 10327 38648 10337 38704
rect 10393 38648 10403 38704
rect 10327 38562 10339 38648
rect 10391 38562 10403 38648
rect 10327 38506 10337 38562
rect 10393 38506 10403 38562
rect 10644 38676 10720 40028
rect 10644 38520 10656 38676
rect 10708 38520 10720 38676
rect 10644 38508 10720 38520
rect 10888 38676 10964 40300
rect 10888 38520 10900 38676
rect 10952 38520 10964 38676
rect 10888 38508 10964 38520
rect 11200 39418 11276 40438
rect 11520 40240 11596 40654
rect 11416 40228 11596 40240
rect 11416 40176 11428 40228
rect 11584 40176 11596 40228
rect 11416 40164 11596 40176
rect 11200 39414 11212 39418
rect 11264 39414 11276 39418
rect 11200 39358 11210 39414
rect 11266 39358 11276 39414
rect 11200 39272 11212 39358
rect 11264 39272 11276 39358
rect 11200 39216 11210 39272
rect 11266 39216 11276 39272
rect 11200 39130 11212 39216
rect 11264 39130 11276 39216
rect 11200 39074 11210 39130
rect 11266 39074 11276 39130
rect 11200 38988 11212 39074
rect 11264 38988 11276 39074
rect 11200 38932 11210 38988
rect 11266 38932 11276 38988
rect 11200 38846 11212 38932
rect 11264 38846 11276 38932
rect 11200 38790 11210 38846
rect 11266 38790 11276 38846
rect 11200 38704 11212 38790
rect 11264 38704 11276 38790
rect 11200 38648 11210 38704
rect 11266 38648 11276 38704
rect 11200 38562 11212 38648
rect 11264 38562 11276 38648
rect 10327 38430 10339 38506
rect 10391 38430 10403 38506
rect 10327 38420 10403 38430
rect 10327 38364 10337 38420
rect 10393 38364 10403 38420
rect 10327 38354 10403 38364
rect 11200 38506 11210 38562
rect 11266 38506 11276 38562
rect 11200 38430 11212 38506
rect 11264 38430 11276 38506
rect 11200 38420 11276 38430
rect 11200 38364 11210 38420
rect 11266 38364 11276 38420
rect 11200 38354 11276 38364
rect 8293 38318 8369 38330
rect 8293 38162 8305 38318
rect 8357 38162 8369 38318
rect 8293 36404 8369 38162
rect 11520 38315 11596 40164
rect 11520 38159 11532 38315
rect 11584 38159 11596 38315
rect 8671 38142 8747 38154
rect 11520 38147 11596 38159
rect 8439 37569 8515 37581
rect 8439 37413 8451 37569
rect 8503 37413 8515 37569
rect 8439 36632 8515 37413
rect 8439 36476 8451 36632
rect 8503 36476 8515 36632
rect 8439 36464 8515 36476
rect 8671 37154 8683 38142
rect 8735 37154 8747 38142
rect 8895 37569 9566 37581
rect 8895 37413 8907 37569
rect 8959 37413 9566 37569
rect 8895 37401 9566 37413
rect 8293 36392 8473 36404
rect 8293 36340 8305 36392
rect 8461 36340 8473 36392
rect 8293 36328 8473 36340
rect 8318 35848 8498 35860
rect 8318 35796 8330 35848
rect 8486 35796 8498 35848
rect 8318 35784 8498 35796
rect 8318 32518 8394 35784
rect 8671 35612 8747 37154
rect 8970 36256 9150 36268
rect 8970 36204 8982 36256
rect 9138 36204 9150 36256
rect 8970 36192 9150 36204
rect 8671 35588 8681 35612
rect 8567 35576 8681 35588
rect 8567 35524 8579 35576
rect 8737 35556 8747 35612
rect 8735 35524 8747 35556
rect 8567 35512 8747 35524
rect 8671 35470 8747 35512
rect 8671 35414 8681 35470
rect 8737 35414 8747 35470
rect 8671 35328 8747 35414
rect 8671 35272 8681 35328
rect 8737 35272 8747 35328
rect 8671 35186 8747 35272
rect 8671 35130 8681 35186
rect 8737 35130 8747 35186
rect 8671 35044 8747 35130
rect 8671 34988 8681 35044
rect 8737 34988 8747 35044
rect 8671 34902 8747 34988
rect 8671 34846 8681 34902
rect 8737 34846 8747 34902
rect 8671 34760 8747 34846
rect 8671 34704 8681 34760
rect 8737 34704 8747 34760
rect 8671 34618 8747 34704
rect 8671 34562 8681 34618
rect 8737 34562 8747 34618
rect 8671 34476 8747 34562
rect 8671 34420 8681 34476
rect 8737 34420 8747 34476
rect 8671 34334 8747 34420
rect 8671 34278 8681 34334
rect 8737 34278 8747 34334
rect 8671 34192 8747 34278
rect 8671 34136 8681 34192
rect 8737 34136 8747 34192
rect 8671 34126 8747 34136
rect 8830 36120 9010 36132
rect 8830 36068 8842 36120
rect 8998 36068 9010 36120
rect 8830 36056 9010 36068
rect 8830 34065 8906 36056
rect 8830 33909 8842 34065
rect 8894 33909 8906 34065
rect 8830 33897 8906 33909
rect 9074 34065 9150 36192
rect 9074 33909 9086 34065
rect 9138 33909 9150 34065
rect 9074 33897 9150 33909
rect 9490 35996 9566 37401
rect 11690 37342 11890 40407
rect 11984 40104 12060 40803
rect 11984 40092 12164 40104
rect 11984 40040 11996 40092
rect 12152 40040 12164 40092
rect 11984 40028 12164 40040
rect 12406 37797 12624 43631
rect 13096 42598 13608 42626
rect 13096 42542 13191 42598
rect 13247 42542 13303 42598
rect 13359 42542 13415 42598
rect 13471 42542 13608 42598
rect 13096 42498 13608 42542
rect 13096 42342 13108 42498
rect 13160 42486 13544 42498
rect 13160 42430 13191 42486
rect 13247 42430 13303 42486
rect 13359 42430 13415 42486
rect 13471 42430 13544 42486
rect 13160 42374 13544 42430
rect 13160 42342 13191 42374
rect 13096 42318 13191 42342
rect 13247 42318 13303 42374
rect 13359 42318 13415 42374
rect 13471 42342 13544 42374
rect 13596 42342 13608 42498
rect 13471 42318 13608 42342
rect 13096 42262 13608 42318
rect 13096 42206 13191 42262
rect 13247 42206 13303 42262
rect 13359 42206 13415 42262
rect 13471 42206 13608 42262
rect 13096 42150 13608 42206
rect 13096 42094 13191 42150
rect 13247 42094 13303 42150
rect 13359 42094 13415 42150
rect 13471 42094 13608 42150
rect 13096 42038 13608 42094
rect 13096 41982 13191 42038
rect 13247 41982 13303 42038
rect 13359 41982 13415 42038
rect 13471 41982 13608 42038
rect 13096 41926 13608 41982
rect 13096 41870 13191 41926
rect 13247 41870 13303 41926
rect 13359 41870 13415 41926
rect 13471 41870 13608 41926
rect 13096 41814 13608 41870
rect 13096 41758 13191 41814
rect 13247 41758 13303 41814
rect 13359 41758 13415 41814
rect 13471 41758 13608 41814
rect 13096 41702 13608 41758
rect 13096 41646 13191 41702
rect 13247 41646 13303 41702
rect 13359 41646 13415 41702
rect 13471 41646 13608 41702
rect 13096 41590 13608 41646
rect 13096 41571 13191 41590
rect 13096 41415 13108 41571
rect 13160 41534 13191 41571
rect 13247 41534 13303 41590
rect 13359 41534 13415 41590
rect 13471 41571 13608 41590
rect 13471 41534 13544 41571
rect 13160 41478 13544 41534
rect 13160 41422 13191 41478
rect 13247 41422 13303 41478
rect 13359 41422 13415 41478
rect 13471 41422 13544 41478
rect 13160 41415 13544 41422
rect 13596 41415 13608 41571
rect 13096 41403 13608 41415
rect 13766 40240 13842 57230
rect 13662 40228 13842 40240
rect 13662 40176 13674 40228
rect 13830 40176 13842 40228
rect 13662 40164 13842 40176
rect 13912 40104 13988 57230
rect 14058 40468 14134 57230
rect 14204 51012 14280 57230
rect 14380 56345 14780 56377
rect 14380 56189 14392 56345
rect 14548 56189 14780 56345
rect 14380 55397 14780 56189
rect 14380 55341 14410 55397
rect 14466 55341 14552 55397
rect 14608 55341 14694 55397
rect 14750 55341 14780 55397
rect 14380 55255 14780 55341
rect 14380 55199 14410 55255
rect 14466 55199 14552 55255
rect 14608 55199 14694 55255
rect 14750 55199 14780 55255
rect 14380 55113 14780 55199
rect 14380 55057 14410 55113
rect 14466 55057 14552 55113
rect 14608 55057 14694 55113
rect 14750 55057 14780 55113
rect 14380 54971 14780 55057
rect 14380 54915 14410 54971
rect 14466 54915 14552 54971
rect 14608 54915 14694 54971
rect 14750 54915 14780 54971
rect 14380 54829 14780 54915
rect 14380 54773 14410 54829
rect 14466 54773 14552 54829
rect 14608 54773 14694 54829
rect 14750 54773 14780 54829
rect 14380 54687 14780 54773
rect 14380 54631 14410 54687
rect 14466 54631 14552 54687
rect 14608 54631 14694 54687
rect 14750 54631 14780 54687
rect 14380 54545 14780 54631
rect 14380 54489 14410 54545
rect 14466 54489 14552 54545
rect 14608 54489 14694 54545
rect 14750 54489 14780 54545
rect 14380 54403 14780 54489
rect 14380 54347 14410 54403
rect 14466 54347 14552 54403
rect 14608 54347 14694 54403
rect 14750 54347 14780 54403
rect 14380 54261 14780 54347
rect 14380 54205 14410 54261
rect 14466 54205 14552 54261
rect 14608 54205 14694 54261
rect 14750 54205 14780 54261
rect 14380 54119 14780 54205
rect 14380 54063 14410 54119
rect 14466 54063 14552 54119
rect 14608 54063 14694 54119
rect 14750 54063 14780 54119
rect 14058 40312 14070 40468
rect 14122 40312 14134 40468
rect 14058 40300 14134 40312
rect 14380 44197 14780 54063
rect 14942 52197 15032 52230
rect 14942 52141 14952 52197
rect 15008 52141 15032 52197
rect 14942 52055 14954 52141
rect 15006 52055 15032 52141
rect 14942 51999 14952 52055
rect 15008 51999 15032 52055
rect 14942 51913 14954 51999
rect 15006 51913 15032 51999
rect 14942 51857 14952 51913
rect 15008 51857 15032 51913
rect 14942 51771 14954 51857
rect 15006 51771 15032 51857
rect 14942 51715 14952 51771
rect 15008 51715 15032 51771
rect 14942 51629 14954 51715
rect 15006 51629 15032 51715
rect 14942 51573 14952 51629
rect 15008 51573 15032 51629
rect 14942 51487 14954 51573
rect 15006 51487 15032 51573
rect 14942 51431 14952 51487
rect 15008 51431 15032 51487
rect 14942 51345 14954 51431
rect 15006 51345 15032 51431
rect 14942 51289 14952 51345
rect 15008 51289 15032 51345
rect 14942 51203 14954 51289
rect 15006 51203 15032 51289
rect 14942 51147 14952 51203
rect 15008 51147 15032 51203
rect 14942 51061 14954 51147
rect 15006 51061 15032 51147
rect 14942 51005 14952 51061
rect 15008 51005 15032 51061
rect 14942 50919 14954 51005
rect 15006 50919 15032 51005
rect 14942 50863 14952 50919
rect 15008 50863 15032 50919
rect 14942 50830 15032 50863
rect 14380 44141 14410 44197
rect 14466 44141 14552 44197
rect 14608 44141 14694 44197
rect 14750 44141 14780 44197
rect 14380 44055 14780 44141
rect 14380 43999 14410 44055
rect 14466 43999 14552 44055
rect 14608 43999 14694 44055
rect 14750 43999 14780 44055
rect 14380 43913 14780 43999
rect 14380 43857 14410 43913
rect 14466 43857 14552 43913
rect 14608 43857 14694 43913
rect 14750 43857 14780 43913
rect 14380 43771 14780 43857
rect 14380 43715 14410 43771
rect 14466 43715 14552 43771
rect 14608 43715 14694 43771
rect 14750 43715 14780 43771
rect 14380 43629 14780 43715
rect 14380 43573 14410 43629
rect 14466 43573 14552 43629
rect 14608 43573 14694 43629
rect 14750 43573 14780 43629
rect 14380 43487 14780 43573
rect 14380 43431 14410 43487
rect 14466 43431 14552 43487
rect 14608 43431 14694 43487
rect 14750 43431 14780 43487
rect 14380 43345 14780 43431
rect 14380 43289 14410 43345
rect 14466 43289 14552 43345
rect 14608 43289 14694 43345
rect 14750 43289 14780 43345
rect 14380 43203 14780 43289
rect 14380 43147 14410 43203
rect 14466 43147 14552 43203
rect 14608 43147 14694 43203
rect 14750 43147 14780 43203
rect 14380 43061 14780 43147
rect 14380 43005 14410 43061
rect 14466 43005 14552 43061
rect 14608 43005 14694 43061
rect 14750 43005 14780 43061
rect 14380 42919 14780 43005
rect 14380 42863 14410 42919
rect 14466 42863 14552 42919
rect 14608 42863 14694 42919
rect 14750 42863 14780 42919
rect 14380 42597 14780 42863
rect 14380 42541 14410 42597
rect 14466 42541 14552 42597
rect 14608 42541 14694 42597
rect 14750 42541 14780 42597
rect 14380 42455 14780 42541
rect 14380 42399 14410 42455
rect 14466 42399 14552 42455
rect 14608 42399 14694 42455
rect 14750 42399 14780 42455
rect 14380 42313 14780 42399
rect 14380 42257 14410 42313
rect 14466 42257 14552 42313
rect 14608 42257 14694 42313
rect 14750 42257 14780 42313
rect 14380 42171 14780 42257
rect 14380 42115 14410 42171
rect 14466 42115 14552 42171
rect 14608 42115 14694 42171
rect 14750 42115 14780 42171
rect 14380 42029 14780 42115
rect 14380 41973 14410 42029
rect 14466 41973 14552 42029
rect 14608 41973 14694 42029
rect 14750 41973 14780 42029
rect 14380 41887 14780 41973
rect 14380 41831 14410 41887
rect 14466 41831 14552 41887
rect 14608 41831 14694 41887
rect 14750 41831 14780 41887
rect 14380 41745 14780 41831
rect 14380 41689 14410 41745
rect 14466 41689 14552 41745
rect 14608 41689 14694 41745
rect 14750 41689 14780 41745
rect 14380 41603 14780 41689
rect 14380 41547 14410 41603
rect 14466 41547 14552 41603
rect 14608 41547 14694 41603
rect 14750 41547 14780 41603
rect 14380 41461 14780 41547
rect 14380 41405 14410 41461
rect 14466 41405 14552 41461
rect 14608 41405 14694 41461
rect 14750 41405 14780 41461
rect 14380 41319 14780 41405
rect 14380 41263 14410 41319
rect 14466 41263 14552 41319
rect 14608 41263 14694 41319
rect 14750 41263 14780 41319
rect 14380 40997 14780 41263
rect 14380 40941 14410 40997
rect 14466 40941 14552 40997
rect 14608 40941 14694 40997
rect 14750 40941 14780 40997
rect 14380 40855 14780 40941
rect 14380 40799 14410 40855
rect 14466 40799 14552 40855
rect 14608 40799 14694 40855
rect 14750 40799 14780 40855
rect 14380 40713 14780 40799
rect 14380 40657 14410 40713
rect 14466 40657 14552 40713
rect 14608 40657 14694 40713
rect 14750 40657 14780 40713
rect 14380 40571 14780 40657
rect 14380 40515 14410 40571
rect 14466 40515 14552 40571
rect 14608 40515 14694 40571
rect 14750 40515 14780 40571
rect 14380 40429 14780 40515
rect 14380 40373 14410 40429
rect 14466 40373 14552 40429
rect 14608 40373 14694 40429
rect 14750 40373 14780 40429
rect 13808 40092 13988 40104
rect 13808 40040 13820 40092
rect 13976 40040 13988 40092
rect 13808 40028 13988 40040
rect 14380 40287 14780 40373
rect 14380 40231 14410 40287
rect 14466 40231 14552 40287
rect 14608 40231 14694 40287
rect 14750 40231 14780 40287
rect 14380 40145 14780 40231
rect 14380 40089 14410 40145
rect 14466 40089 14552 40145
rect 14608 40089 14694 40145
rect 14750 40089 14780 40145
rect 14380 40003 14780 40089
rect 12748 39946 13818 39956
rect 12748 39890 12758 39946
rect 12814 39944 12900 39946
rect 12956 39944 13042 39946
rect 13098 39944 13184 39946
rect 13240 39944 13326 39946
rect 13382 39944 13468 39946
rect 13524 39944 13610 39946
rect 13666 39944 13752 39946
rect 12814 39890 12900 39892
rect 12956 39890 13042 39892
rect 13098 39890 13184 39892
rect 13240 39890 13326 39892
rect 13382 39890 13468 39892
rect 13524 39890 13610 39892
rect 13666 39890 13752 39892
rect 13808 39890 13818 39946
rect 12748 39880 13818 39890
rect 14380 39947 14410 40003
rect 14466 39947 14552 40003
rect 14608 39947 14694 40003
rect 14750 39947 14780 40003
rect 14380 39861 14780 39947
rect 14380 39805 14410 39861
rect 14466 39805 14552 39861
rect 14608 39805 14694 39861
rect 14750 39805 14780 39861
rect 14380 39719 14780 39805
rect 14380 39663 14410 39719
rect 14466 39663 14552 39719
rect 14608 39663 14694 39719
rect 14750 39663 14780 39719
rect 13303 38307 13754 38319
rect 13303 38151 13315 38307
rect 13367 38151 13754 38307
rect 13303 38139 13754 38151
rect 12406 37741 12416 37797
rect 12472 37741 12558 37797
rect 12614 37741 12624 37797
rect 12406 37655 12624 37741
rect 12406 37599 12416 37655
rect 12472 37599 12558 37655
rect 12614 37599 12624 37655
rect 12406 37513 12624 37599
rect 12406 37457 12416 37513
rect 12472 37457 12558 37513
rect 12614 37457 12624 37513
rect 12406 37371 12624 37457
rect 10331 37200 11551 37210
rect 10331 37198 10435 37200
rect 10491 37198 10577 37200
rect 10633 37198 10719 37200
rect 10775 37198 10861 37200
rect 10917 37198 11003 37200
rect 11059 37198 11145 37200
rect 11201 37198 11287 37200
rect 11343 37198 11429 37200
rect 11485 37198 11551 37200
rect 10331 37146 10343 37198
rect 11539 37146 11551 37198
rect 10331 37144 10435 37146
rect 10491 37144 10577 37146
rect 10633 37144 10719 37146
rect 10775 37144 10861 37146
rect 10917 37144 11003 37146
rect 11059 37144 11145 37146
rect 11201 37144 11287 37146
rect 11343 37144 11429 37146
rect 11485 37144 11551 37146
rect 10331 37134 11551 37144
rect 11690 37142 12090 37342
rect 9490 35984 9670 35996
rect 9490 35932 9502 35984
rect 9658 35932 9670 35984
rect 9490 35920 9670 35932
rect 9490 34065 9566 35920
rect 10394 35712 10574 35724
rect 10394 35660 10406 35712
rect 10562 35660 10574 35712
rect 10394 35648 10574 35660
rect 10998 35716 11074 35726
rect 10998 35660 11008 35716
rect 11064 35660 11074 35716
rect 10100 35612 10176 35622
rect 10100 35556 10110 35612
rect 10166 35556 10176 35612
rect 10100 35470 10112 35556
rect 10164 35470 10176 35556
rect 10100 35414 10110 35470
rect 10166 35414 10176 35470
rect 10100 35328 10112 35414
rect 10164 35328 10176 35414
rect 10100 35272 10110 35328
rect 10166 35272 10176 35328
rect 10100 35186 10112 35272
rect 10164 35186 10176 35272
rect 10100 35130 10110 35186
rect 10166 35130 10176 35186
rect 10100 35044 10112 35130
rect 10164 35044 10176 35130
rect 10100 34988 10110 35044
rect 10166 34988 10176 35044
rect 10100 34902 10112 34988
rect 10164 34902 10176 34988
rect 10100 34846 10110 34902
rect 10166 34846 10176 34902
rect 10100 34760 10112 34846
rect 10164 34760 10176 34846
rect 10100 34704 10110 34760
rect 10166 34704 10176 34760
rect 10100 34618 10112 34704
rect 10164 34618 10176 34704
rect 10100 34562 10110 34618
rect 10166 34562 10176 34618
rect 10100 34476 10112 34562
rect 10164 34476 10176 34562
rect 10100 34420 10110 34476
rect 10166 34420 10176 34476
rect 10100 34334 10112 34420
rect 10164 34334 10176 34420
rect 10100 34278 10110 34334
rect 10166 34278 10176 34334
rect 10100 34192 10112 34278
rect 10164 34192 10176 34278
rect 10100 34136 10110 34192
rect 10166 34136 10176 34192
rect 10100 34126 10176 34136
rect 9490 33909 9502 34065
rect 9554 33909 9566 34065
rect 9490 33897 9566 33909
rect 10394 33897 10470 35648
rect 10998 35576 11074 35660
rect 11498 35712 11678 35724
rect 11498 35660 11510 35712
rect 11666 35660 11678 35712
rect 11498 35648 11678 35660
rect 10998 35574 11010 35576
rect 11062 35574 11074 35576
rect 10998 35518 11008 35574
rect 11064 35518 11074 35574
rect 10998 35432 11010 35518
rect 11062 35432 11074 35518
rect 10998 35376 11008 35432
rect 11064 35376 11074 35432
rect 10998 35290 11010 35376
rect 11062 35290 11074 35376
rect 10998 35234 11008 35290
rect 11064 35234 11074 35290
rect 10998 35148 11010 35234
rect 11062 35148 11074 35234
rect 10998 35092 11008 35148
rect 11064 35092 11074 35148
rect 10998 35006 11010 35092
rect 11062 35006 11074 35092
rect 10998 34950 11008 35006
rect 11064 34950 11074 35006
rect 10998 34864 11010 34950
rect 11062 34864 11074 34950
rect 10998 34808 11008 34864
rect 11064 34808 11074 34864
rect 10998 34722 11010 34808
rect 11062 34722 11074 34808
rect 10998 34666 11008 34722
rect 11064 34666 11074 34722
rect 10998 34580 11010 34666
rect 11062 34580 11074 34666
rect 10998 34524 11008 34580
rect 11064 34524 11074 34580
rect 10998 34438 11010 34524
rect 11062 34438 11074 34524
rect 10998 34382 11008 34438
rect 11064 34382 11074 34438
rect 10998 34296 11010 34382
rect 11062 34296 11074 34382
rect 10998 34240 11008 34296
rect 11064 34240 11074 34296
rect 10998 34154 11010 34240
rect 11062 34154 11074 34240
rect 10998 34098 11008 34154
rect 11064 34098 11074 34154
rect 10998 34012 11010 34098
rect 11062 34012 11074 34098
rect 10998 33956 11008 34012
rect 11064 33956 11074 34012
rect 10998 33870 11010 33956
rect 11062 33870 11074 33956
rect 11602 33897 11678 35648
rect 11890 35612 12090 37142
rect 12406 37315 12416 37371
rect 12472 37315 12558 37371
rect 12614 37315 12624 37371
rect 12406 37229 12624 37315
rect 12406 37173 12416 37229
rect 12472 37173 12558 37229
rect 12614 37173 12624 37229
rect 12406 37087 12624 37173
rect 12406 37031 12416 37087
rect 12472 37031 12558 37087
rect 12614 37031 12624 37087
rect 12406 36945 12624 37031
rect 12406 36889 12416 36945
rect 12472 36889 12558 36945
rect 12614 36889 12624 36945
rect 12406 36803 12624 36889
rect 12406 36747 12416 36803
rect 12472 36747 12558 36803
rect 12614 36747 12624 36803
rect 12406 36661 12624 36747
rect 12406 36605 12416 36661
rect 12472 36605 12558 36661
rect 12614 36605 12624 36661
rect 12406 36519 12624 36605
rect 13439 37653 13515 37665
rect 13439 37497 13451 37653
rect 13503 37497 13515 37653
rect 12406 36463 12416 36519
rect 12472 36463 12558 36519
rect 12614 36463 12624 36519
rect 13062 36528 13242 36540
rect 13062 36476 13074 36528
rect 13230 36476 13242 36528
rect 13062 36464 13242 36476
rect 12406 36430 12624 36463
rect 12922 36392 13102 36404
rect 12922 36340 12934 36392
rect 13090 36340 13102 36392
rect 12922 36328 13102 36340
rect 11890 35556 11906 35612
rect 11962 35556 12090 35612
rect 11890 35470 11908 35556
rect 11960 35470 12090 35556
rect 11890 35414 11906 35470
rect 11962 35414 12090 35470
rect 11890 35328 11908 35414
rect 11960 35328 12090 35414
rect 11890 35272 11906 35328
rect 11962 35272 12090 35328
rect 11890 35186 11908 35272
rect 11960 35186 12090 35272
rect 11890 35130 11906 35186
rect 11962 35130 12090 35186
rect 11890 35044 11908 35130
rect 11960 35044 12090 35130
rect 11890 34988 11906 35044
rect 11962 34988 12090 35044
rect 11890 34902 11908 34988
rect 11960 34902 12090 34988
rect 11890 34846 11906 34902
rect 11962 34846 12090 34902
rect 11890 34760 11908 34846
rect 11960 34760 12090 34846
rect 11890 34704 11906 34760
rect 11962 34704 12090 34760
rect 11890 34618 11908 34704
rect 11960 34618 12090 34704
rect 11890 34562 11906 34618
rect 11962 34562 12090 34618
rect 11890 34476 11908 34562
rect 11960 34476 12090 34562
rect 11890 34420 11906 34476
rect 11962 34420 12090 34476
rect 11890 34334 11908 34420
rect 11960 34334 12090 34420
rect 11890 34278 11906 34334
rect 11962 34278 12090 34334
rect 11890 34192 11908 34278
rect 11960 34192 12090 34278
rect 11890 34136 11906 34192
rect 11962 34136 12090 34192
rect 11890 34129 12090 34136
rect 12506 35984 12686 35996
rect 12506 35932 12518 35984
rect 12674 35932 12686 35984
rect 12506 35920 12686 35932
rect 11896 34126 11972 34129
rect 12506 34065 12582 35920
rect 12506 33909 12518 34065
rect 12570 33909 12582 34065
rect 12506 33897 12582 33909
rect 12922 34065 12998 36328
rect 12922 33909 12934 34065
rect 12986 33909 12998 34065
rect 12922 33897 12998 33909
rect 13166 34065 13242 36464
rect 13439 35724 13515 37497
rect 13678 35860 13754 38139
rect 13574 35848 13754 35860
rect 13574 35796 13586 35848
rect 13742 35796 13754 35848
rect 13574 35784 13754 35796
rect 13335 35712 13515 35724
rect 13335 35660 13347 35712
rect 13503 35660 13515 35712
rect 13335 35648 13515 35660
rect 13166 33909 13178 34065
rect 13230 33909 13242 34065
rect 13166 33897 13242 33909
rect 10998 33814 11008 33870
rect 11064 33814 11074 33870
rect 10998 33728 11010 33814
rect 11062 33728 11074 33814
rect 10998 33672 11008 33728
rect 11064 33672 11074 33728
rect 10998 33586 11010 33672
rect 11062 33586 11074 33672
rect 10998 33530 11008 33586
rect 11064 33530 11074 33586
rect 10998 33444 11010 33530
rect 11062 33444 11074 33530
rect 10998 33388 11008 33444
rect 11064 33388 11074 33444
rect 10998 33302 11010 33388
rect 11062 33302 11074 33388
rect 10998 33246 11008 33302
rect 11064 33246 11074 33302
rect 10998 32924 11010 33246
rect 11062 32924 11074 33246
rect 10998 32912 11074 32924
rect 10998 32535 11074 32545
rect 10998 32479 11008 32535
rect 11064 32479 11074 32535
rect 13678 32518 13754 35784
rect 14380 33481 14780 39663
rect 14942 37797 15032 37830
rect 14942 37741 14952 37797
rect 15008 37741 15032 37797
rect 14942 37655 14954 37741
rect 15006 37655 15032 37741
rect 14942 37599 14952 37655
rect 15008 37599 15032 37655
rect 14942 37513 14954 37599
rect 15006 37513 15032 37599
rect 14942 37457 14952 37513
rect 15008 37457 15032 37513
rect 14942 37371 14954 37457
rect 15006 37371 15032 37457
rect 14942 37315 14952 37371
rect 15008 37315 15032 37371
rect 14942 37229 14954 37315
rect 15006 37229 15032 37315
rect 14942 37173 14952 37229
rect 15008 37173 15032 37229
rect 14942 37087 14954 37173
rect 15006 37087 15032 37173
rect 14942 37031 14952 37087
rect 15008 37031 15032 37087
rect 14942 36945 14954 37031
rect 15006 36945 15032 37031
rect 14942 36889 14952 36945
rect 15008 36889 15032 36945
rect 14942 36803 14954 36889
rect 15006 36803 15032 36889
rect 14942 36747 14952 36803
rect 15008 36747 15032 36803
rect 14942 36661 14954 36747
rect 15006 36661 15032 36747
rect 14942 36605 14952 36661
rect 15008 36605 15032 36661
rect 14942 36519 14954 36605
rect 15006 36519 15032 36605
rect 14942 36463 14952 36519
rect 15008 36463 15032 36519
rect 14942 36430 15032 36463
rect 14380 32978 14514 33481
rect 14566 32978 14780 33481
rect 14380 32922 14410 32978
rect 14466 32922 14514 32978
rect 14608 32922 14694 32978
rect 14750 32922 14780 32978
rect 14380 32836 14514 32922
rect 14566 32836 14780 32922
rect 14380 32780 14410 32836
rect 14466 32780 14514 32836
rect 14608 32780 14694 32836
rect 14750 32780 14780 32836
rect 14380 32694 14514 32780
rect 14566 32694 14780 32780
rect 14380 32638 14410 32694
rect 14466 32638 14514 32694
rect 14608 32638 14694 32694
rect 14750 32638 14780 32694
rect 14380 32552 14514 32638
rect 14566 32552 14780 32638
rect 10998 32455 11074 32479
rect 10998 32393 11010 32455
rect 11062 32393 11074 32455
rect 10998 32337 11008 32393
rect 11064 32337 11074 32393
rect 7976 32322 8052 32332
rect 7976 32266 7986 32322
rect 8042 32266 8052 32322
rect 7976 32180 7988 32266
rect 8040 32180 8052 32266
rect 7976 32124 7986 32180
rect 8042 32124 8052 32180
rect 7976 32038 7988 32124
rect 8040 32038 8052 32124
rect 7976 31982 7986 32038
rect 8042 31982 8052 32038
rect 7976 31896 7988 31982
rect 8040 31896 8052 31982
rect 7976 31840 7986 31896
rect 8042 31840 8052 31896
rect 7976 31754 7988 31840
rect 8040 31754 8052 31840
rect 7976 31698 7986 31754
rect 8042 31698 8052 31754
rect 7976 31612 7988 31698
rect 8040 31612 8052 31698
rect 7976 31556 7986 31612
rect 8042 31556 8052 31612
rect 7976 31470 7988 31556
rect 8040 31470 8052 31556
rect 7976 31414 7986 31470
rect 8042 31414 8052 31470
rect 7976 31328 7988 31414
rect 8040 31328 8052 31414
rect 7976 31272 7986 31328
rect 8042 31272 8052 31328
rect 7976 31186 7988 31272
rect 8040 31186 8052 31272
rect 7976 31130 7986 31186
rect 8042 31130 8052 31186
rect 7976 31044 7988 31130
rect 8040 31044 8052 31130
rect 7976 30988 7986 31044
rect 8042 30988 8052 31044
rect 7976 30902 7988 30988
rect 8040 30902 8052 30988
rect 7976 30846 7986 30902
rect 8042 30846 8052 30902
rect 7976 30760 7988 30846
rect 8040 30760 8052 30846
rect 7976 30704 7986 30760
rect 8042 30704 8052 30760
rect 7976 30618 7988 30704
rect 8040 30618 8052 30704
rect 9368 32323 9444 32333
rect 9368 32267 9378 32323
rect 9434 32267 9444 32323
rect 9368 32181 9380 32267
rect 9432 32181 9444 32267
rect 9368 32125 9378 32181
rect 9434 32125 9444 32181
rect 9368 32039 9380 32125
rect 9432 32039 9444 32125
rect 9368 31983 9378 32039
rect 9434 31983 9444 32039
rect 9368 31897 9380 31983
rect 9432 31897 9444 31983
rect 9368 31841 9378 31897
rect 9434 31841 9444 31897
rect 9368 31755 9380 31841
rect 9432 31755 9444 31841
rect 9368 31699 9378 31755
rect 9434 31699 9444 31755
rect 9368 31613 9380 31699
rect 9432 31613 9444 31699
rect 9368 31557 9378 31613
rect 9434 31557 9444 31613
rect 9368 31471 9380 31557
rect 9432 31471 9444 31557
rect 9368 31415 9378 31471
rect 9434 31415 9444 31471
rect 9368 31329 9380 31415
rect 9432 31329 9444 31415
rect 9368 31273 9378 31329
rect 9434 31273 9444 31329
rect 9368 31187 9380 31273
rect 9432 31187 9444 31273
rect 9368 31131 9378 31187
rect 9434 31131 9444 31187
rect 9368 31045 9380 31131
rect 9432 31045 9444 31131
rect 9368 30989 9378 31045
rect 9434 30989 9444 31045
rect 9368 30903 9380 30989
rect 9432 30903 9444 30989
rect 9368 30847 9378 30903
rect 9434 30847 9444 30903
rect 9368 30761 9380 30847
rect 9432 30761 9444 30847
rect 9368 30705 9378 30761
rect 9434 30705 9444 30761
rect 9368 30695 9444 30705
rect 9784 32323 9860 32333
rect 9784 32267 9794 32323
rect 9850 32267 9860 32323
rect 9784 32181 9796 32267
rect 9848 32181 9860 32267
rect 9784 32125 9794 32181
rect 9850 32125 9860 32181
rect 9784 32039 9796 32125
rect 9848 32039 9860 32125
rect 9784 31983 9794 32039
rect 9850 31983 9860 32039
rect 9784 31897 9796 31983
rect 9848 31897 9860 31983
rect 9784 31841 9794 31897
rect 9850 31841 9860 31897
rect 9784 31755 9796 31841
rect 9848 31755 9860 31841
rect 9784 31699 9794 31755
rect 9850 31699 9860 31755
rect 9784 31613 9796 31699
rect 9848 31613 9860 31699
rect 9784 31557 9794 31613
rect 9850 31557 9860 31613
rect 9784 31471 9796 31557
rect 9848 31471 9860 31557
rect 9784 31415 9794 31471
rect 9850 31415 9860 31471
rect 9784 31329 9796 31415
rect 9848 31329 9860 31415
rect 9784 31273 9794 31329
rect 9850 31273 9860 31329
rect 9784 31187 9796 31273
rect 9848 31187 9860 31273
rect 9784 31131 9794 31187
rect 9850 31131 9860 31187
rect 9784 31045 9796 31131
rect 9848 31045 9860 31131
rect 9784 30989 9794 31045
rect 9850 30989 9860 31045
rect 9784 30903 9796 30989
rect 9848 30903 9860 30989
rect 9784 30847 9794 30903
rect 9850 30847 9860 30903
rect 9784 30761 9796 30847
rect 9848 30761 9860 30847
rect 9784 30705 9794 30761
rect 9850 30705 9860 30761
rect 9784 30695 9860 30705
rect 10272 32323 10348 32333
rect 10272 32267 10282 32323
rect 10338 32267 10348 32323
rect 10272 32181 10284 32267
rect 10336 32181 10348 32267
rect 10272 32125 10282 32181
rect 10338 32125 10348 32181
rect 10272 32039 10284 32125
rect 10336 32039 10348 32125
rect 10272 31983 10282 32039
rect 10338 31983 10348 32039
rect 10272 31897 10284 31983
rect 10336 31897 10348 31983
rect 10272 31841 10282 31897
rect 10338 31841 10348 31897
rect 10272 31755 10284 31841
rect 10336 31755 10348 31841
rect 10272 31699 10282 31755
rect 10338 31699 10348 31755
rect 10272 31613 10284 31699
rect 10336 31613 10348 31699
rect 10272 31557 10282 31613
rect 10338 31557 10348 31613
rect 10272 31471 10284 31557
rect 10336 31471 10348 31557
rect 10272 31415 10282 31471
rect 10338 31415 10348 31471
rect 10272 31329 10284 31415
rect 10336 31329 10348 31415
rect 10272 31273 10282 31329
rect 10338 31273 10348 31329
rect 10272 31187 10284 31273
rect 10336 31187 10348 31273
rect 10272 31131 10282 31187
rect 10338 31131 10348 31187
rect 10272 31045 10284 31131
rect 10336 31045 10348 31131
rect 10272 30989 10282 31045
rect 10338 30989 10348 31045
rect 10272 30903 10284 30989
rect 10336 30903 10348 30989
rect 10272 30847 10282 30903
rect 10338 30847 10348 30903
rect 10272 30761 10284 30847
rect 10336 30761 10348 30847
rect 10272 30705 10282 30761
rect 10338 30705 10348 30761
rect 10272 30695 10348 30705
rect 10760 32272 10836 32282
rect 10760 32216 10770 32272
rect 10826 32216 10836 32272
rect 10760 32130 10772 32216
rect 10824 32130 10836 32216
rect 10760 32074 10770 32130
rect 10826 32074 10836 32130
rect 10760 31988 10772 32074
rect 10824 31988 10836 32074
rect 10760 31932 10770 31988
rect 10826 31932 10836 31988
rect 10760 31846 10772 31932
rect 10824 31846 10836 31932
rect 10760 31790 10770 31846
rect 10826 31790 10836 31846
rect 10760 31704 10772 31790
rect 10824 31704 10836 31790
rect 10760 31648 10770 31704
rect 10826 31648 10836 31704
rect 10760 31562 10772 31648
rect 10824 31562 10836 31648
rect 10760 31506 10770 31562
rect 10826 31506 10836 31562
rect 10760 31420 10772 31506
rect 10824 31420 10836 31506
rect 10760 31364 10770 31420
rect 10826 31364 10836 31420
rect 10760 31278 10772 31364
rect 10824 31278 10836 31364
rect 10760 31222 10770 31278
rect 10826 31222 10836 31278
rect 10760 31136 10772 31222
rect 10824 31136 10836 31222
rect 10760 31080 10770 31136
rect 10826 31080 10836 31136
rect 10760 30994 10772 31080
rect 10824 30994 10836 31080
rect 10760 30938 10770 30994
rect 10826 30938 10836 30994
rect 10760 30852 10772 30938
rect 10824 30852 10836 30938
rect 10760 30796 10770 30852
rect 10826 30796 10836 30852
rect 10760 30710 10772 30796
rect 10824 30710 10836 30796
rect 10760 30654 10770 30710
rect 10826 30654 10836 30710
rect 10760 30644 10836 30654
rect 10998 32251 11010 32337
rect 11062 32251 11074 32337
rect 14380 32496 14410 32552
rect 14466 32496 14514 32552
rect 14608 32496 14694 32552
rect 14750 32496 14780 32552
rect 14380 32410 14514 32496
rect 14566 32410 14780 32496
rect 14380 32354 14410 32410
rect 14466 32354 14514 32410
rect 14608 32354 14694 32410
rect 14750 32354 14780 32410
rect 11724 32323 11800 32333
rect 10998 32195 11008 32251
rect 11064 32195 11074 32251
rect 10998 32109 11010 32195
rect 11062 32109 11074 32195
rect 10998 32053 11008 32109
rect 11064 32053 11074 32109
rect 10998 31967 11010 32053
rect 11062 31967 11074 32053
rect 10998 31911 11008 31967
rect 11064 31911 11074 31967
rect 10998 31825 11010 31911
rect 11062 31825 11074 31911
rect 10998 31769 11008 31825
rect 11064 31769 11074 31825
rect 10998 31683 11010 31769
rect 11062 31683 11074 31769
rect 10998 31627 11008 31683
rect 11064 31627 11074 31683
rect 10998 31541 11010 31627
rect 11062 31541 11074 31627
rect 10998 31485 11008 31541
rect 11064 31485 11074 31541
rect 10998 31399 11010 31485
rect 11062 31399 11074 31485
rect 10998 31343 11008 31399
rect 11064 31343 11074 31399
rect 10998 31257 11010 31343
rect 11062 31257 11074 31343
rect 10998 31201 11008 31257
rect 11064 31201 11074 31257
rect 10998 31115 11010 31201
rect 11062 31115 11074 31201
rect 10998 31059 11008 31115
rect 11064 31059 11074 31115
rect 10998 30973 11010 31059
rect 11062 30973 11074 31059
rect 10998 30917 11008 30973
rect 11064 30917 11074 30973
rect 10998 30831 11010 30917
rect 11062 30831 11074 30917
rect 10998 30775 11008 30831
rect 11064 30775 11074 30831
rect 10998 30689 11010 30775
rect 11062 30689 11074 30775
rect 10998 30633 11008 30689
rect 11064 30633 11074 30689
rect 11236 32272 11312 32282
rect 11236 32216 11246 32272
rect 11302 32216 11312 32272
rect 11236 32130 11248 32216
rect 11300 32130 11312 32216
rect 11236 32074 11246 32130
rect 11302 32074 11312 32130
rect 11236 31988 11248 32074
rect 11300 31988 11312 32074
rect 11236 31932 11246 31988
rect 11302 31932 11312 31988
rect 11236 31846 11248 31932
rect 11300 31846 11312 31932
rect 11236 31790 11246 31846
rect 11302 31790 11312 31846
rect 11236 31704 11248 31790
rect 11300 31704 11312 31790
rect 11236 31648 11246 31704
rect 11302 31648 11312 31704
rect 11236 31562 11248 31648
rect 11300 31562 11312 31648
rect 11236 31506 11246 31562
rect 11302 31506 11312 31562
rect 11236 31420 11248 31506
rect 11300 31420 11312 31506
rect 11236 31364 11246 31420
rect 11302 31364 11312 31420
rect 11236 31278 11248 31364
rect 11300 31278 11312 31364
rect 11236 31222 11246 31278
rect 11302 31222 11312 31278
rect 11236 31136 11248 31222
rect 11300 31136 11312 31222
rect 11236 31080 11246 31136
rect 11302 31080 11312 31136
rect 11236 30994 11248 31080
rect 11300 30994 11312 31080
rect 11236 30938 11246 30994
rect 11302 30938 11312 30994
rect 11236 30852 11248 30938
rect 11300 30852 11312 30938
rect 11236 30796 11246 30852
rect 11302 30796 11312 30852
rect 11236 30710 11248 30796
rect 11300 30710 11312 30796
rect 11236 30654 11246 30710
rect 11302 30654 11312 30710
rect 11724 32267 11734 32323
rect 11790 32267 11800 32323
rect 11724 32181 11736 32267
rect 11788 32181 11800 32267
rect 11724 32125 11734 32181
rect 11790 32125 11800 32181
rect 11724 32039 11736 32125
rect 11788 32039 11800 32125
rect 11724 31983 11734 32039
rect 11790 31983 11800 32039
rect 11724 31897 11736 31983
rect 11788 31897 11800 31983
rect 11724 31841 11734 31897
rect 11790 31841 11800 31897
rect 11724 31755 11736 31841
rect 11788 31755 11800 31841
rect 11724 31699 11734 31755
rect 11790 31699 11800 31755
rect 11724 31613 11736 31699
rect 11788 31613 11800 31699
rect 11724 31557 11734 31613
rect 11790 31557 11800 31613
rect 11724 31471 11736 31557
rect 11788 31471 11800 31557
rect 11724 31415 11734 31471
rect 11790 31415 11800 31471
rect 11724 31329 11736 31415
rect 11788 31329 11800 31415
rect 11724 31273 11734 31329
rect 11790 31273 11800 31329
rect 11724 31187 11736 31273
rect 11788 31187 11800 31273
rect 11724 31131 11734 31187
rect 11790 31131 11800 31187
rect 11724 31045 11736 31131
rect 11788 31045 11800 31131
rect 11724 30989 11734 31045
rect 11790 30989 11800 31045
rect 11724 30903 11736 30989
rect 11788 30903 11800 30989
rect 11724 30847 11734 30903
rect 11790 30847 11800 30903
rect 11724 30761 11736 30847
rect 11788 30761 11800 30847
rect 11724 30705 11734 30761
rect 11790 30705 11800 30761
rect 11724 30695 11800 30705
rect 12212 32322 12288 32332
rect 12212 32266 12222 32322
rect 12278 32266 12288 32322
rect 12212 32180 12224 32266
rect 12276 32180 12288 32266
rect 12212 32124 12222 32180
rect 12278 32124 12288 32180
rect 12212 32038 12224 32124
rect 12276 32038 12288 32124
rect 12212 31982 12222 32038
rect 12278 31982 12288 32038
rect 12212 31896 12224 31982
rect 12276 31896 12288 31982
rect 12212 31840 12222 31896
rect 12278 31840 12288 31896
rect 12212 31754 12224 31840
rect 12276 31754 12288 31840
rect 12212 31698 12222 31754
rect 12278 31698 12288 31754
rect 12212 31612 12224 31698
rect 12276 31612 12288 31698
rect 12212 31556 12222 31612
rect 12278 31556 12288 31612
rect 12212 31470 12224 31556
rect 12276 31470 12288 31556
rect 12212 31414 12222 31470
rect 12278 31414 12288 31470
rect 12212 31328 12224 31414
rect 12276 31328 12288 31414
rect 12212 31272 12222 31328
rect 12278 31272 12288 31328
rect 12212 31186 12224 31272
rect 12276 31186 12288 31272
rect 12212 31130 12222 31186
rect 12278 31130 12288 31186
rect 12212 31044 12224 31130
rect 12276 31044 12288 31130
rect 12212 30988 12222 31044
rect 12278 30988 12288 31044
rect 12212 30902 12224 30988
rect 12276 30902 12288 30988
rect 12212 30846 12222 30902
rect 12278 30846 12288 30902
rect 12212 30760 12224 30846
rect 12276 30760 12288 30846
rect 12212 30704 12222 30760
rect 12278 30704 12288 30760
rect 11236 30644 11312 30654
rect 10998 30623 11074 30633
rect 7976 30562 7986 30618
rect 8042 30562 8052 30618
rect 7976 30476 7988 30562
rect 8040 30476 8052 30562
rect 12212 30618 12224 30704
rect 12276 30618 12288 30704
rect 12212 30562 12222 30618
rect 12278 30562 12288 30618
rect 7976 30420 7986 30476
rect 8042 30420 8052 30476
rect 7976 30334 7988 30420
rect 8040 30334 8052 30420
rect 7976 30278 7986 30334
rect 8042 30278 8052 30334
rect 9062 30488 10592 30500
rect 9062 30400 10528 30488
rect 7976 30192 7988 30278
rect 8040 30192 8052 30278
rect 7976 30136 7986 30192
rect 8042 30136 8052 30192
rect 7976 30084 7988 30136
rect 8040 30084 8052 30136
rect 7976 30072 8052 30084
rect 8452 30308 8552 30320
rect 8452 29944 8476 30308
rect 8528 29944 8552 30308
rect 8452 29279 8552 29944
rect 8696 30308 8796 30320
rect 8696 29944 8720 30308
rect 8772 29944 8796 30308
rect 8696 29459 8796 29944
rect 8696 29447 8876 29459
rect 8696 29395 8708 29447
rect 8864 29395 8876 29447
rect 8696 29383 8876 29395
rect 8452 29267 8632 29279
rect 8452 29215 8464 29267
rect 8620 29215 8632 29267
rect 8452 29203 8632 29215
rect 9062 29099 9162 30400
rect 9062 28943 9088 29099
rect 9140 28943 9162 29099
rect 9062 28931 9162 28943
rect 10016 30308 10116 30320
rect 10016 29944 10040 30308
rect 10092 29944 10116 30308
rect 10516 30124 10528 30400
rect 10580 30124 10592 30488
rect 10516 30112 10592 30124
rect 10821 30488 12044 30500
rect 10821 30400 11980 30488
rect 10016 29099 10116 29944
rect 10016 28943 10042 29099
rect 10094 28943 10116 29099
rect 10016 28931 10116 28943
rect 10821 29099 10921 30400
rect 10821 28943 10847 29099
rect 10899 28943 10921 29099
rect 11468 30308 11568 30320
rect 11468 29944 11492 30308
rect 11544 29944 11568 30308
rect 11968 30124 11980 30400
rect 12032 30124 12044 30488
rect 11968 30112 12044 30124
rect 12212 30476 12224 30562
rect 12276 30476 12288 30562
rect 12212 30420 12222 30476
rect 12278 30420 12288 30476
rect 12212 30334 12224 30420
rect 12276 30334 12288 30420
rect 12212 30278 12222 30334
rect 12278 30278 12288 30334
rect 12212 30192 12224 30278
rect 12276 30192 12288 30278
rect 12212 30136 12222 30192
rect 12278 30136 12288 30192
rect 12212 30084 12224 30136
rect 12276 30084 12288 30136
rect 12212 30072 12288 30084
rect 12628 32322 12704 32332
rect 12628 32266 12638 32322
rect 12694 32266 12704 32322
rect 12628 32180 12640 32266
rect 12692 32180 12704 32266
rect 12628 32124 12638 32180
rect 12694 32124 12704 32180
rect 12628 32038 12640 32124
rect 12692 32038 12704 32124
rect 12628 31982 12638 32038
rect 12694 31982 12704 32038
rect 12628 31896 12640 31982
rect 12692 31896 12704 31982
rect 12628 31840 12638 31896
rect 12694 31840 12704 31896
rect 12628 31754 12640 31840
rect 12692 31754 12704 31840
rect 12628 31698 12638 31754
rect 12694 31698 12704 31754
rect 12628 31612 12640 31698
rect 12692 31612 12704 31698
rect 12628 31556 12638 31612
rect 12694 31556 12704 31612
rect 12628 31470 12640 31556
rect 12692 31470 12704 31556
rect 12628 31414 12638 31470
rect 12694 31414 12704 31470
rect 12628 31328 12640 31414
rect 12692 31328 12704 31414
rect 12628 31272 12638 31328
rect 12694 31272 12704 31328
rect 12628 31186 12640 31272
rect 12692 31186 12704 31272
rect 12628 31130 12638 31186
rect 12694 31130 12704 31186
rect 12628 31044 12640 31130
rect 12692 31044 12704 31130
rect 12628 30988 12638 31044
rect 12694 30988 12704 31044
rect 12628 30902 12640 30988
rect 12692 30902 12704 30988
rect 12628 30846 12638 30902
rect 12694 30846 12704 30902
rect 12628 30760 12640 30846
rect 12692 30760 12704 30846
rect 12628 30704 12638 30760
rect 12694 30704 12704 30760
rect 12628 30618 12640 30704
rect 12692 30618 12704 30704
rect 12628 30562 12638 30618
rect 12694 30562 12704 30618
rect 12628 30476 12640 30562
rect 12692 30476 12704 30562
rect 12628 30420 12638 30476
rect 12694 30420 12704 30476
rect 12628 30334 12640 30420
rect 12692 30334 12704 30420
rect 12628 30278 12638 30334
rect 12694 30278 12704 30334
rect 14020 32322 14096 32332
rect 14020 32266 14030 32322
rect 14086 32266 14096 32322
rect 14020 32180 14032 32266
rect 14084 32180 14096 32266
rect 14020 32124 14030 32180
rect 14086 32124 14096 32180
rect 14020 32038 14032 32124
rect 14084 32038 14096 32124
rect 14020 31982 14030 32038
rect 14086 31982 14096 32038
rect 14020 31896 14032 31982
rect 14084 31896 14096 31982
rect 14020 31840 14030 31896
rect 14086 31840 14096 31896
rect 14020 31754 14032 31840
rect 14084 31754 14096 31840
rect 14020 31698 14030 31754
rect 14086 31698 14096 31754
rect 14020 31612 14032 31698
rect 14084 31612 14096 31698
rect 14020 31556 14030 31612
rect 14086 31556 14096 31612
rect 14020 31470 14032 31556
rect 14084 31470 14096 31556
rect 14020 31414 14030 31470
rect 14086 31414 14096 31470
rect 14020 31328 14032 31414
rect 14084 31328 14096 31414
rect 14020 31272 14030 31328
rect 14086 31272 14096 31328
rect 14020 31186 14032 31272
rect 14084 31186 14096 31272
rect 14020 31130 14030 31186
rect 14086 31130 14096 31186
rect 14020 31044 14032 31130
rect 14084 31044 14096 31130
rect 14020 30988 14030 31044
rect 14086 30988 14096 31044
rect 14020 30902 14032 30988
rect 14084 30902 14096 30988
rect 14020 30846 14030 30902
rect 14086 30846 14096 30902
rect 14020 30760 14032 30846
rect 14084 30760 14096 30846
rect 14020 30704 14030 30760
rect 14086 30704 14096 30760
rect 14020 30618 14032 30704
rect 14084 30618 14096 30704
rect 14020 30562 14030 30618
rect 14086 30562 14096 30618
rect 14020 30476 14032 30562
rect 14084 30476 14096 30562
rect 14020 30420 14030 30476
rect 14086 30420 14096 30476
rect 14020 30334 14032 30420
rect 14084 30334 14096 30420
rect 12628 30192 12640 30278
rect 12692 30192 12704 30278
rect 12628 30136 12638 30192
rect 12694 30136 12704 30192
rect 12628 30084 12640 30136
rect 12692 30084 12704 30136
rect 12628 30072 12704 30084
rect 13520 30308 13620 30320
rect 11468 29072 11568 29944
rect 13520 29944 13544 30308
rect 13596 29944 13620 30308
rect 11922 29739 13276 29749
rect 11922 29683 11932 29739
rect 11988 29737 12074 29739
rect 12130 29737 12216 29739
rect 12272 29737 12358 29739
rect 12414 29737 12500 29739
rect 12556 29737 12642 29739
rect 12698 29737 12784 29739
rect 12840 29737 12926 29739
rect 12982 29737 13068 29739
rect 13124 29737 13210 29739
rect 11988 29683 12074 29685
rect 12130 29683 12216 29685
rect 12272 29683 12358 29685
rect 12414 29683 12500 29685
rect 12556 29683 12642 29685
rect 12698 29683 12784 29685
rect 12840 29683 12926 29685
rect 12982 29683 13068 29685
rect 13124 29683 13210 29685
rect 13266 29683 13276 29739
rect 11922 29673 13276 29683
rect 13520 29651 13620 29944
rect 13764 30308 13864 30320
rect 13764 29944 13788 30308
rect 13840 29944 13864 30308
rect 14020 30278 14030 30334
rect 14086 30278 14096 30334
rect 14020 30192 14032 30278
rect 14084 30192 14096 30278
rect 14020 30136 14030 30192
rect 14086 30136 14096 30192
rect 14020 30084 14032 30136
rect 14084 30084 14096 30136
rect 14020 30072 14096 30084
rect 14380 32268 14514 32354
rect 14566 32268 14780 32354
rect 14380 32212 14410 32268
rect 14466 32212 14514 32268
rect 14608 32212 14694 32268
rect 14750 32212 14780 32268
rect 14380 32126 14514 32212
rect 14566 32126 14780 32212
rect 14380 32070 14410 32126
rect 14466 32070 14514 32126
rect 14608 32070 14694 32126
rect 14750 32070 14780 32126
rect 14380 31984 14514 32070
rect 14566 31984 14780 32070
rect 14380 31928 14410 31984
rect 14466 31928 14514 31984
rect 14608 31928 14694 31984
rect 14750 31928 14780 31984
rect 14380 31842 14514 31928
rect 14566 31842 14780 31928
rect 14380 31786 14410 31842
rect 14466 31786 14514 31842
rect 14608 31786 14694 31842
rect 14750 31786 14780 31842
rect 14380 31700 14514 31786
rect 14566 31700 14780 31786
rect 14380 31644 14410 31700
rect 14466 31644 14514 31700
rect 14608 31644 14694 31700
rect 14750 31644 14780 31700
rect 14380 31558 14514 31644
rect 14566 31558 14780 31644
rect 14380 31502 14410 31558
rect 14466 31502 14514 31558
rect 14608 31502 14694 31558
rect 14750 31502 14780 31558
rect 14380 31416 14514 31502
rect 14566 31416 14780 31502
rect 14380 31360 14410 31416
rect 14466 31360 14514 31416
rect 14608 31360 14694 31416
rect 14750 31360 14780 31416
rect 14380 31274 14514 31360
rect 14566 31274 14780 31360
rect 14380 31218 14410 31274
rect 14466 31218 14514 31274
rect 14608 31218 14694 31274
rect 14750 31218 14780 31274
rect 14380 31132 14514 31218
rect 14566 31132 14780 31218
rect 14380 31076 14410 31132
rect 14466 31076 14514 31132
rect 14608 31076 14694 31132
rect 14750 31076 14780 31132
rect 14380 30990 14514 31076
rect 14566 30990 14780 31076
rect 14380 30934 14410 30990
rect 14466 30934 14514 30990
rect 14608 30934 14694 30990
rect 14750 30934 14780 30990
rect 14380 30848 14514 30934
rect 14566 30848 14780 30934
rect 14380 30792 14410 30848
rect 14466 30792 14514 30848
rect 14608 30792 14694 30848
rect 14750 30792 14780 30848
rect 14380 30706 14514 30792
rect 14566 30706 14780 30792
rect 14380 30650 14410 30706
rect 14466 30650 14514 30706
rect 14608 30650 14694 30706
rect 14750 30650 14780 30706
rect 14380 30564 14514 30650
rect 14566 30564 14780 30650
rect 14380 30508 14410 30564
rect 14466 30508 14514 30564
rect 14608 30508 14694 30564
rect 14750 30508 14780 30564
rect 14380 30422 14514 30508
rect 14566 30422 14780 30508
rect 14380 30366 14410 30422
rect 14466 30366 14514 30422
rect 14608 30366 14694 30422
rect 14750 30366 14780 30422
rect 14380 30280 14514 30366
rect 14566 30280 14780 30366
rect 14380 30224 14410 30280
rect 14466 30224 14514 30280
rect 14608 30224 14694 30280
rect 14750 30224 14780 30280
rect 14380 30138 14514 30224
rect 14566 30138 14780 30224
rect 14380 30082 14410 30138
rect 14466 30082 14514 30138
rect 14608 30082 14694 30138
rect 14750 30082 14780 30138
rect 13764 29831 13864 29944
rect 13764 29731 14059 29831
rect 13520 29551 13879 29651
rect 13519 29447 13699 29459
rect 13519 29395 13531 29447
rect 13687 29395 13699 29447
rect 13519 29383 13699 29395
rect 13339 29267 13519 29279
rect 13339 29215 13351 29267
rect 13507 29215 13519 29267
rect 13339 29203 13519 29215
rect 11390 29060 11570 29072
rect 11390 29008 11402 29060
rect 11558 29008 11570 29060
rect 11390 28996 11570 29008
rect 10821 28931 10921 28943
rect 13411 28031 13519 29203
rect 13599 28031 13699 29383
rect 13779 28031 13879 29551
rect 13959 28031 14059 29731
rect 14380 29797 14514 30082
rect 14566 29797 14780 30082
rect 14380 29741 14410 29797
rect 14466 29741 14514 29797
rect 14608 29741 14694 29797
rect 14750 29741 14780 29797
rect 14380 29685 14514 29741
rect 14566 29685 14780 29741
rect 14380 29655 14780 29685
rect 14380 29599 14410 29655
rect 14466 29599 14552 29655
rect 14608 29599 14694 29655
rect 14750 29599 14780 29655
rect 14380 29513 14780 29599
rect 14380 29457 14410 29513
rect 14466 29457 14552 29513
rect 14608 29457 14694 29513
rect 14750 29457 14780 29513
rect 14380 29371 14780 29457
rect 14380 29315 14410 29371
rect 14466 29315 14552 29371
rect 14608 29315 14694 29371
rect 14750 29315 14780 29371
rect 14380 29229 14780 29315
rect 14380 29173 14410 29229
rect 14466 29173 14552 29229
rect 14608 29173 14694 29229
rect 14750 29173 14780 29229
rect 14380 29087 14780 29173
rect 14380 29031 14410 29087
rect 14466 29031 14552 29087
rect 14608 29031 14694 29087
rect 14750 29031 14780 29087
rect 14380 28945 14780 29031
rect 14380 28889 14410 28945
rect 14466 28889 14552 28945
rect 14608 28889 14694 28945
rect 14750 28889 14780 28945
rect 14380 28803 14780 28889
rect 14380 28747 14410 28803
rect 14466 28747 14552 28803
rect 14608 28747 14694 28803
rect 14750 28747 14780 28803
rect 14380 28661 14780 28747
rect 14380 28605 14410 28661
rect 14466 28605 14552 28661
rect 14608 28605 14694 28661
rect 14750 28605 14780 28661
rect 14380 28519 14780 28605
rect 14380 28463 14410 28519
rect 14466 28463 14552 28519
rect 14608 28463 14694 28519
rect 14750 28463 14780 28519
rect 165 27573 175 27629
rect 231 27573 317 27629
rect 373 27573 383 27629
rect 165 27487 383 27573
rect 165 27431 175 27487
rect 231 27431 317 27487
rect 373 27431 383 27487
rect 165 27345 383 27431
rect 165 27289 175 27345
rect 231 27289 317 27345
rect 373 27289 383 27345
rect 165 27203 383 27289
rect 165 27147 175 27203
rect 231 27147 317 27203
rect 373 27147 383 27203
rect 165 27061 383 27147
rect 165 27005 175 27061
rect 231 27005 317 27061
rect 373 27005 383 27061
rect 165 26919 383 27005
rect 165 26863 175 26919
rect 231 26863 317 26919
rect 373 26863 383 26919
rect 165 13744 383 26863
rect 14380 26578 14780 28463
rect 14380 26522 14410 26578
rect 14466 26522 14552 26578
rect 14608 26522 14694 26578
rect 14750 26522 14780 26578
rect 14380 26436 14780 26522
rect 14380 26380 14410 26436
rect 14466 26380 14552 26436
rect 14608 26380 14694 26436
rect 14750 26380 14780 26436
rect 14380 26294 14780 26380
rect 14380 26238 14410 26294
rect 14466 26238 14552 26294
rect 14608 26238 14694 26294
rect 14750 26238 14780 26294
rect 14380 26152 14780 26238
rect 14380 26096 14410 26152
rect 14466 26096 14552 26152
rect 14608 26096 14694 26152
rect 14750 26096 14780 26152
rect 14380 26010 14780 26096
rect 14380 25954 14410 26010
rect 14466 25954 14552 26010
rect 14608 25954 14694 26010
rect 14750 25954 14780 26010
rect 14380 25868 14780 25954
rect 14380 25812 14410 25868
rect 14466 25812 14552 25868
rect 14608 25812 14694 25868
rect 14750 25812 14780 25868
rect 14380 25726 14780 25812
rect 14380 25670 14410 25726
rect 14466 25670 14552 25726
rect 14608 25670 14694 25726
rect 14750 25670 14780 25726
rect 14380 25584 14780 25670
rect 14380 25528 14410 25584
rect 14466 25528 14552 25584
rect 14608 25528 14694 25584
rect 14750 25528 14780 25584
rect 14380 25442 14780 25528
rect 14380 25386 14410 25442
rect 14466 25386 14552 25442
rect 14608 25386 14694 25442
rect 14750 25386 14780 25442
rect 14380 25300 14780 25386
rect 14380 25244 14410 25300
rect 14466 25244 14552 25300
rect 14608 25244 14694 25300
rect 14750 25244 14780 25300
rect 14380 25158 14780 25244
rect 14380 25102 14410 25158
rect 14466 25102 14552 25158
rect 14608 25102 14694 25158
rect 14750 25102 14780 25158
rect 14380 25016 14780 25102
rect 14380 24960 14410 25016
rect 14466 24960 14552 25016
rect 14608 24960 14694 25016
rect 14750 24960 14780 25016
rect 14380 24874 14780 24960
rect 14380 24818 14410 24874
rect 14466 24818 14552 24874
rect 14608 24818 14694 24874
rect 14750 24818 14780 24874
rect 14380 24732 14780 24818
rect 14380 24676 14410 24732
rect 14466 24676 14552 24732
rect 14608 24676 14694 24732
rect 14750 24676 14780 24732
rect 14380 24590 14780 24676
rect 14380 24534 14410 24590
rect 14466 24534 14552 24590
rect 14608 24534 14694 24590
rect 14750 24534 14780 24590
rect 14380 24448 14780 24534
rect 14380 24392 14410 24448
rect 14466 24392 14552 24448
rect 14608 24392 14694 24448
rect 14750 24392 14780 24448
rect 14380 24306 14780 24392
rect 14380 24250 14410 24306
rect 14466 24250 14552 24306
rect 14608 24250 14694 24306
rect 14750 24250 14780 24306
rect 14380 24164 14780 24250
rect 14380 24108 14410 24164
rect 14466 24108 14552 24164
rect 14608 24108 14694 24164
rect 14750 24108 14780 24164
rect 14380 24022 14780 24108
rect 14380 23966 14410 24022
rect 14466 23966 14552 24022
rect 14608 23966 14694 24022
rect 14750 23966 14780 24022
rect 14380 23880 14780 23966
rect 14380 23824 14410 23880
rect 14466 23824 14552 23880
rect 14608 23824 14694 23880
rect 14750 23824 14780 23880
rect 14380 23738 14780 23824
rect 14380 23682 14410 23738
rect 14466 23682 14552 23738
rect 14608 23682 14694 23738
rect 14750 23682 14780 23738
rect 14380 23378 14780 23682
rect 14380 23322 14410 23378
rect 14466 23322 14552 23378
rect 14608 23322 14694 23378
rect 14750 23322 14780 23378
rect 14380 23236 14780 23322
rect 14380 23180 14410 23236
rect 14466 23180 14552 23236
rect 14608 23180 14694 23236
rect 14750 23180 14780 23236
rect 14380 23094 14780 23180
rect 14380 23038 14410 23094
rect 14466 23038 14552 23094
rect 14608 23038 14694 23094
rect 14750 23038 14780 23094
rect 14380 22952 14780 23038
rect 14380 22896 14410 22952
rect 14466 22896 14552 22952
rect 14608 22896 14694 22952
rect 14750 22896 14780 22952
rect 14380 22810 14780 22896
rect 14380 22754 14410 22810
rect 14466 22754 14552 22810
rect 14608 22754 14694 22810
rect 14750 22754 14780 22810
rect 14380 22668 14780 22754
rect 14380 22612 14410 22668
rect 14466 22612 14552 22668
rect 14608 22612 14694 22668
rect 14750 22612 14780 22668
rect 14380 22526 14780 22612
rect 14380 22470 14410 22526
rect 14466 22470 14552 22526
rect 14608 22470 14694 22526
rect 14750 22470 14780 22526
rect 14380 22384 14780 22470
rect 14380 22328 14410 22384
rect 14466 22328 14552 22384
rect 14608 22328 14694 22384
rect 14750 22328 14780 22384
rect 14380 22242 14780 22328
rect 14380 22186 14410 22242
rect 14466 22186 14552 22242
rect 14608 22186 14694 22242
rect 14750 22186 14780 22242
rect 14380 22100 14780 22186
rect 14380 22044 14410 22100
rect 14466 22044 14552 22100
rect 14608 22044 14694 22100
rect 14750 22044 14780 22100
rect 14380 21958 14780 22044
rect 14380 21902 14410 21958
rect 14466 21902 14552 21958
rect 14608 21902 14694 21958
rect 14750 21902 14780 21958
rect 14380 21816 14780 21902
rect 14380 21760 14410 21816
rect 14466 21760 14552 21816
rect 14608 21760 14694 21816
rect 14750 21760 14780 21816
rect 14380 21674 14780 21760
rect 14380 21618 14410 21674
rect 14466 21618 14552 21674
rect 14608 21618 14694 21674
rect 14750 21618 14780 21674
rect 14380 21532 14780 21618
rect 14380 21476 14410 21532
rect 14466 21476 14552 21532
rect 14608 21476 14694 21532
rect 14750 21476 14780 21532
rect 14380 21390 14780 21476
rect 14380 21334 14410 21390
rect 14466 21334 14552 21390
rect 14608 21334 14694 21390
rect 14750 21334 14780 21390
rect 14380 21248 14780 21334
rect 14380 21192 14410 21248
rect 14466 21192 14552 21248
rect 14608 21192 14694 21248
rect 14750 21192 14780 21248
rect 14380 21106 14780 21192
rect 14380 21050 14410 21106
rect 14466 21050 14552 21106
rect 14608 21050 14694 21106
rect 14750 21050 14780 21106
rect 14380 20964 14780 21050
rect 14380 20908 14410 20964
rect 14466 20908 14552 20964
rect 14608 20908 14694 20964
rect 14750 20908 14780 20964
rect 14380 20822 14780 20908
rect 14380 20766 14410 20822
rect 14466 20766 14552 20822
rect 14608 20766 14694 20822
rect 14750 20766 14780 20822
rect 14380 20680 14780 20766
rect 14380 20624 14410 20680
rect 14466 20624 14552 20680
rect 14608 20624 14694 20680
rect 14750 20624 14780 20680
rect 14380 20538 14780 20624
rect 14380 20482 14410 20538
rect 14466 20482 14552 20538
rect 14608 20482 14694 20538
rect 14750 20482 14780 20538
rect 14380 20178 14780 20482
rect 14380 20122 14410 20178
rect 14466 20122 14552 20178
rect 14608 20122 14694 20178
rect 14750 20122 14780 20178
rect 14380 20036 14780 20122
rect 14380 19980 14410 20036
rect 14466 19980 14552 20036
rect 14608 19980 14694 20036
rect 14750 19980 14780 20036
rect 14380 19894 14780 19980
rect 14380 19838 14410 19894
rect 14466 19838 14552 19894
rect 14608 19838 14694 19894
rect 14750 19838 14780 19894
rect 14380 19752 14780 19838
rect 14380 19696 14410 19752
rect 14466 19696 14552 19752
rect 14608 19696 14694 19752
rect 14750 19696 14780 19752
rect 14380 19610 14780 19696
rect 14380 19554 14410 19610
rect 14466 19554 14552 19610
rect 14608 19554 14694 19610
rect 14750 19554 14780 19610
rect 14380 19468 14780 19554
rect 14380 19412 14410 19468
rect 14466 19412 14552 19468
rect 14608 19412 14694 19468
rect 14750 19412 14780 19468
rect 14380 19326 14780 19412
rect 14380 19270 14410 19326
rect 14466 19270 14552 19326
rect 14608 19270 14694 19326
rect 14750 19270 14780 19326
rect 14380 19184 14780 19270
rect 14380 19128 14410 19184
rect 14466 19128 14552 19184
rect 14608 19128 14694 19184
rect 14750 19128 14780 19184
rect 14380 19042 14780 19128
rect 14380 18986 14410 19042
rect 14466 18986 14552 19042
rect 14608 18986 14694 19042
rect 14750 18986 14780 19042
rect 14380 18900 14780 18986
rect 14380 18844 14410 18900
rect 14466 18844 14552 18900
rect 14608 18844 14694 18900
rect 14750 18844 14780 18900
rect 14380 18758 14780 18844
rect 14380 18702 14410 18758
rect 14466 18702 14552 18758
rect 14608 18702 14694 18758
rect 14750 18702 14780 18758
rect 14380 18616 14780 18702
rect 14380 18560 14410 18616
rect 14466 18560 14552 18616
rect 14608 18560 14694 18616
rect 14750 18560 14780 18616
rect 14380 18474 14780 18560
rect 14380 18418 14410 18474
rect 14466 18418 14552 18474
rect 14608 18418 14694 18474
rect 14750 18418 14780 18474
rect 14380 18332 14780 18418
rect 14380 18276 14410 18332
rect 14466 18276 14552 18332
rect 14608 18276 14694 18332
rect 14750 18276 14780 18332
rect 14380 18190 14780 18276
rect 14380 18134 14410 18190
rect 14466 18134 14552 18190
rect 14608 18134 14694 18190
rect 14750 18134 14780 18190
rect 14380 18048 14780 18134
rect 14380 17992 14410 18048
rect 14466 17992 14552 18048
rect 14608 17992 14694 18048
rect 14750 17992 14780 18048
rect 14380 17906 14780 17992
rect 14380 17850 14410 17906
rect 14466 17850 14552 17906
rect 14608 17850 14694 17906
rect 14750 17850 14780 17906
rect 14380 17764 14780 17850
rect 14380 17708 14410 17764
rect 14466 17708 14552 17764
rect 14608 17708 14694 17764
rect 14750 17708 14780 17764
rect 14380 17622 14780 17708
rect 14380 17566 14410 17622
rect 14466 17566 14552 17622
rect 14608 17566 14694 17622
rect 14750 17566 14780 17622
rect 14380 17480 14780 17566
rect 14380 17424 14410 17480
rect 14466 17424 14552 17480
rect 14608 17424 14694 17480
rect 14750 17424 14780 17480
rect 14380 17338 14780 17424
rect 14380 17282 14410 17338
rect 14466 17282 14552 17338
rect 14608 17282 14694 17338
rect 14750 17282 14780 17338
rect 14380 17030 14780 17282
rect 14380 16978 14834 17030
rect 14380 16922 14410 16978
rect 14466 16922 14552 16978
rect 14608 16922 14694 16978
rect 14750 16922 14834 16978
rect 14380 16836 14834 16922
rect 14380 16780 14410 16836
rect 14466 16780 14552 16836
rect 14608 16780 14694 16836
rect 14750 16780 14834 16836
rect 14380 16694 14834 16780
rect 14380 16638 14410 16694
rect 14466 16638 14552 16694
rect 14608 16638 14694 16694
rect 14750 16638 14834 16694
rect 14380 16552 14834 16638
rect 14380 16496 14410 16552
rect 14466 16496 14552 16552
rect 14608 16496 14694 16552
rect 14750 16496 14834 16552
rect 14380 16410 14834 16496
rect 14380 16354 14410 16410
rect 14466 16354 14552 16410
rect 14608 16354 14694 16410
rect 14750 16354 14834 16410
rect 14380 16268 14834 16354
rect 14380 16212 14410 16268
rect 14466 16212 14552 16268
rect 14608 16212 14694 16268
rect 14750 16212 14834 16268
rect 14380 16126 14834 16212
rect 14380 16070 14410 16126
rect 14466 16070 14552 16126
rect 14608 16070 14694 16126
rect 14750 16070 14834 16126
rect 14380 15984 14834 16070
rect 14380 15928 14410 15984
rect 14466 15928 14552 15984
rect 14608 15928 14694 15984
rect 14750 15928 14834 15984
rect 14380 15842 14834 15928
rect 14380 15786 14410 15842
rect 14466 15786 14552 15842
rect 14608 15786 14694 15842
rect 14750 15786 14834 15842
rect 14380 15700 14834 15786
rect 14380 15644 14410 15700
rect 14466 15644 14552 15700
rect 14608 15644 14694 15700
rect 14750 15644 14834 15700
rect 14380 15558 14834 15644
rect 14380 15502 14410 15558
rect 14466 15502 14552 15558
rect 14608 15502 14694 15558
rect 14750 15502 14834 15558
rect 14380 15416 14834 15502
rect 14380 15360 14410 15416
rect 14466 15360 14552 15416
rect 14608 15360 14694 15416
rect 14750 15360 14834 15416
rect 14380 15274 14834 15360
rect 14380 15218 14410 15274
rect 14466 15218 14552 15274
rect 14608 15218 14694 15274
rect 14750 15218 14834 15274
rect 14380 15132 14834 15218
rect 14380 15076 14410 15132
rect 14466 15076 14552 15132
rect 14608 15076 14694 15132
rect 14750 15076 14834 15132
rect 14380 14990 14834 15076
rect 14380 14934 14410 14990
rect 14466 14934 14552 14990
rect 14608 14934 14694 14990
rect 14750 14934 14834 14990
rect 14380 14848 14834 14934
rect 14380 14792 14410 14848
rect 14466 14792 14552 14848
rect 14608 14792 14694 14848
rect 14750 14792 14834 14848
rect 14380 14706 14834 14792
rect 14380 14650 14410 14706
rect 14466 14650 14552 14706
rect 14608 14650 14694 14706
rect 14750 14650 14834 14706
rect 14380 14564 14834 14650
rect 14380 14508 14410 14564
rect 14466 14508 14552 14564
rect 14608 14508 14694 14564
rect 14750 14508 14834 14564
rect 14380 14422 14834 14508
rect 14380 14366 14410 14422
rect 14466 14366 14552 14422
rect 14608 14366 14694 14422
rect 14750 14366 14834 14422
rect 14380 14280 14834 14366
rect 14380 14224 14410 14280
rect 14466 14224 14552 14280
rect 14608 14224 14694 14280
rect 14750 14224 14834 14280
rect 14380 14138 14834 14224
rect 14380 14082 14410 14138
rect 14466 14082 14552 14138
rect 14608 14082 14694 14138
rect 14750 14082 14834 14138
rect 14380 14030 14834 14082
rect 165 12524 870 13744
rect 165 10578 383 12524
rect 14634 11923 14834 14030
rect 14169 10853 14834 11923
rect 165 10522 175 10578
rect 231 10522 317 10578
rect 373 10522 383 10578
rect 165 10436 383 10522
rect 165 10380 175 10436
rect 231 10380 317 10436
rect 373 10380 383 10436
rect 165 10294 383 10380
rect 165 10238 175 10294
rect 231 10238 317 10294
rect 373 10238 383 10294
rect 165 10152 383 10238
rect 165 10096 175 10152
rect 231 10096 317 10152
rect 373 10096 383 10152
rect 165 10010 383 10096
rect 165 9954 175 10010
rect 231 9954 317 10010
rect 373 9954 383 10010
rect 165 9868 383 9954
rect 165 9812 175 9868
rect 231 9812 317 9868
rect 373 9812 383 9868
rect 165 9726 383 9812
rect 165 9670 175 9726
rect 231 9670 317 9726
rect 373 9670 383 9726
rect 165 9584 383 9670
rect 165 9528 175 9584
rect 231 9528 317 9584
rect 373 9528 383 9584
rect 165 9442 383 9528
rect 165 9386 175 9442
rect 231 9386 317 9442
rect 373 9386 383 9442
rect 165 9300 383 9386
rect 165 9244 175 9300
rect 231 9244 317 9300
rect 373 9244 383 9300
rect 165 9158 383 9244
rect 165 9102 175 9158
rect 231 9102 317 9158
rect 373 9102 383 9158
rect 165 9016 383 9102
rect 165 8960 175 9016
rect 231 8960 317 9016
rect 373 8960 383 9016
rect 165 8874 383 8960
rect 165 8818 175 8874
rect 231 8818 317 8874
rect 373 8818 383 8874
rect 165 8732 383 8818
rect 165 8676 175 8732
rect 231 8676 317 8732
rect 373 8676 383 8732
rect 165 8590 383 8676
rect 165 8534 175 8590
rect 231 8534 317 8590
rect 373 8534 383 8590
rect 165 8448 383 8534
rect 165 8392 175 8448
rect 231 8392 317 8448
rect 373 8392 383 8448
rect 165 8306 383 8392
rect 165 8250 175 8306
rect 231 8250 317 8306
rect 373 8250 383 8306
rect 165 8164 383 8250
rect 165 8108 175 8164
rect 231 8108 317 8164
rect 373 8108 383 8164
rect 165 8022 383 8108
rect 165 7966 175 8022
rect 231 7966 317 8022
rect 373 7966 383 8022
rect 165 7880 383 7966
rect 165 7824 175 7880
rect 231 7824 317 7880
rect 373 7824 383 7880
rect 165 7738 383 7824
rect 165 7682 175 7738
rect 231 7682 317 7738
rect 373 7682 383 7738
rect 165 7378 383 7682
rect 165 7322 175 7378
rect 231 7322 317 7378
rect 373 7322 383 7378
rect 165 7236 383 7322
rect 165 7180 175 7236
rect 231 7180 317 7236
rect 373 7180 383 7236
rect 165 7094 383 7180
rect 165 7038 175 7094
rect 231 7038 317 7094
rect 373 7038 383 7094
rect 165 6952 383 7038
rect 165 6896 175 6952
rect 231 6896 317 6952
rect 373 6896 383 6952
rect 165 6810 383 6896
rect 165 6754 175 6810
rect 231 6754 317 6810
rect 373 6754 383 6810
rect 165 6668 383 6754
rect 165 6612 175 6668
rect 231 6612 317 6668
rect 373 6612 383 6668
rect 165 6526 383 6612
rect 165 6470 175 6526
rect 231 6470 317 6526
rect 373 6470 383 6526
rect 165 6384 383 6470
rect 165 6328 175 6384
rect 231 6328 317 6384
rect 373 6328 383 6384
rect 165 6242 383 6328
rect 165 6186 175 6242
rect 231 6186 317 6242
rect 373 6186 383 6242
rect 165 6100 383 6186
rect 165 6044 175 6100
rect 231 6044 317 6100
rect 373 6044 383 6100
rect 165 5958 383 6044
rect 165 5902 175 5958
rect 231 5902 317 5958
rect 373 5902 383 5958
rect 165 5816 383 5902
rect 165 5760 175 5816
rect 231 5760 317 5816
rect 373 5760 383 5816
rect 165 5674 383 5760
rect 165 5618 175 5674
rect 231 5618 317 5674
rect 373 5618 383 5674
rect 165 5532 383 5618
rect 165 5476 175 5532
rect 231 5476 317 5532
rect 373 5476 383 5532
rect 165 5390 383 5476
rect 165 5334 175 5390
rect 231 5334 317 5390
rect 373 5334 383 5390
rect 165 5248 383 5334
rect 165 5192 175 5248
rect 231 5192 317 5248
rect 373 5192 383 5248
rect 165 5106 383 5192
rect 165 5050 175 5106
rect 231 5050 317 5106
rect 373 5050 383 5106
rect 165 4964 383 5050
rect 165 4908 175 4964
rect 231 4908 317 4964
rect 373 4908 383 4964
rect 165 4822 383 4908
rect 165 4766 175 4822
rect 231 4766 317 4822
rect 373 4766 383 4822
rect 165 4680 383 4766
rect 165 4624 175 4680
rect 231 4624 317 4680
rect 373 4624 383 4680
rect 165 4538 383 4624
rect 165 4482 175 4538
rect 231 4482 317 4538
rect 373 4482 383 4538
rect 165 4178 383 4482
rect 165 4122 175 4178
rect 231 4122 317 4178
rect 373 4122 383 4178
rect 165 4036 383 4122
rect 165 3980 175 4036
rect 231 3980 317 4036
rect 373 3980 383 4036
rect 165 3894 383 3980
rect 165 3838 175 3894
rect 231 3838 317 3894
rect 373 3838 383 3894
rect 165 3752 383 3838
rect 165 3696 175 3752
rect 231 3696 317 3752
rect 373 3696 383 3752
rect 165 3610 383 3696
rect 165 3554 175 3610
rect 231 3554 317 3610
rect 373 3554 383 3610
rect 165 3468 383 3554
rect 165 3412 175 3468
rect 231 3412 317 3468
rect 373 3412 383 3468
rect 165 3326 383 3412
rect 165 3270 175 3326
rect 231 3270 317 3326
rect 373 3270 383 3326
rect 165 3184 383 3270
rect 165 3128 175 3184
rect 231 3128 317 3184
rect 373 3128 383 3184
rect 165 3042 383 3128
rect 165 2986 175 3042
rect 231 2986 317 3042
rect 373 2986 383 3042
rect 165 2900 383 2986
rect 165 2844 175 2900
rect 231 2844 317 2900
rect 373 2844 383 2900
rect 165 2758 383 2844
rect 165 2702 175 2758
rect 231 2702 317 2758
rect 373 2702 383 2758
rect 165 2616 383 2702
rect 165 2560 175 2616
rect 231 2560 317 2616
rect 373 2560 383 2616
rect 165 2474 383 2560
rect 165 2418 175 2474
rect 231 2418 317 2474
rect 373 2418 383 2474
rect 165 2332 383 2418
rect 165 2276 175 2332
rect 231 2276 317 2332
rect 373 2276 383 2332
rect 165 2190 383 2276
rect 165 2134 175 2190
rect 231 2134 317 2190
rect 373 2134 383 2190
rect 165 2048 383 2134
rect 165 1992 175 2048
rect 231 1992 317 2048
rect 373 1992 383 2048
rect 165 1906 383 1992
rect 165 1850 175 1906
rect 231 1850 317 1906
rect 373 1850 383 1906
rect 165 1764 383 1850
rect 165 1708 175 1764
rect 231 1708 317 1764
rect 373 1708 383 1764
rect 165 1622 383 1708
rect 165 1566 175 1622
rect 231 1566 317 1622
rect 373 1566 383 1622
rect 165 1480 383 1566
rect 165 1424 175 1480
rect 231 1424 317 1480
rect 373 1424 383 1480
rect 165 1338 383 1424
rect 165 1282 175 1338
rect 231 1282 317 1338
rect 373 1282 383 1338
rect 165 1230 383 1282
<< via2 >>
rect 1896 56809 1952 56865
rect 1896 56667 1952 56723
rect 1896 56525 1952 56581
rect 1896 56383 1952 56439
rect 1896 56241 1952 56297
rect 1896 56099 1952 56155
rect 1896 55957 1952 56013
rect 1896 55815 1952 55871
rect 1896 55673 1952 55729
rect 56 52180 112 52197
rect 56 52141 58 52180
rect 58 52141 110 52180
rect 110 52141 112 52180
rect 56 51999 58 52055
rect 58 51999 110 52055
rect 110 51999 112 52055
rect 56 51857 58 51913
rect 58 51857 110 51913
rect 110 51857 112 51913
rect 56 51715 58 51771
rect 58 51715 110 51771
rect 110 51715 112 51771
rect 56 51573 58 51629
rect 58 51573 110 51629
rect 110 51573 112 51629
rect 56 51431 58 51487
rect 58 51431 110 51487
rect 110 51431 112 51487
rect 56 51289 58 51345
rect 58 51289 110 51345
rect 110 51289 112 51345
rect 56 51147 58 51203
rect 58 51147 110 51203
rect 110 51147 112 51203
rect 56 51005 58 51061
rect 58 51005 110 51061
rect 110 51005 112 51061
rect 56 50880 58 50919
rect 58 50880 110 50919
rect 110 50880 112 50919
rect 56 50863 112 50880
rect 214 50541 270 50597
rect 356 50541 412 50597
rect 498 50541 554 50597
rect 214 50399 270 50455
rect 356 50399 412 50455
rect 498 50399 554 50455
rect 214 50257 270 50313
rect 356 50257 412 50313
rect 498 50257 554 50313
rect 214 50115 270 50171
rect 356 50115 412 50171
rect 498 50115 554 50171
rect 214 49973 270 50029
rect 356 49973 412 50029
rect 498 49973 554 50029
rect 214 49831 270 49887
rect 356 49831 412 49887
rect 498 49831 554 49887
rect 214 49689 270 49745
rect 356 49689 412 49745
rect 498 49689 554 49745
rect 214 49547 270 49603
rect 356 49547 412 49603
rect 498 49547 554 49603
rect 214 49405 270 49461
rect 356 49405 412 49461
rect 498 49405 554 49461
rect 214 49263 270 49319
rect 356 49263 412 49319
rect 498 49263 554 49319
rect 214 39341 270 39397
rect 356 39341 412 39397
rect 498 39341 554 39397
rect 214 39199 270 39255
rect 356 39199 412 39255
rect 498 39199 554 39255
rect 214 39057 270 39113
rect 356 39057 412 39113
rect 498 39057 554 39113
rect 214 38915 270 38971
rect 356 38915 412 38971
rect 498 38915 554 38971
rect 214 38773 270 38829
rect 356 38773 412 38829
rect 498 38773 554 38829
rect 214 38631 270 38687
rect 356 38631 412 38687
rect 498 38631 554 38687
rect 214 38489 270 38545
rect 356 38489 412 38545
rect 498 38489 554 38545
rect 214 38347 270 38403
rect 356 38347 412 38403
rect 498 38347 554 38403
rect 214 38205 270 38261
rect 356 38205 412 38261
rect 498 38205 554 38261
rect 214 38063 270 38119
rect 356 38063 412 38119
rect 498 38063 554 38119
rect 734 52141 790 52197
rect 876 52141 932 52197
rect 1018 52141 1074 52197
rect 734 51999 790 52055
rect 876 51999 932 52055
rect 1018 51999 1074 52055
rect 734 51857 790 51913
rect 876 51857 932 51913
rect 1018 51857 1074 51913
rect 734 51715 790 51771
rect 876 51715 932 51771
rect 1018 51715 1074 51771
rect 734 51573 790 51629
rect 876 51573 932 51629
rect 1018 51573 1074 51629
rect 734 51431 790 51487
rect 876 51431 932 51487
rect 1018 51431 1074 51487
rect 734 51289 790 51345
rect 876 51289 932 51345
rect 1018 51289 1074 51345
rect 734 51147 790 51203
rect 876 51147 932 51203
rect 1018 51147 1074 51203
rect 734 51005 790 51061
rect 876 51005 932 51061
rect 1018 51005 1074 51061
rect 734 50863 790 50919
rect 876 50863 932 50919
rect 1018 50863 1074 50919
rect 1896 53741 1952 53797
rect 1896 53599 1952 53655
rect 1896 53457 1952 53513
rect 1896 53315 1952 53371
rect 1896 53173 1952 53229
rect 2500 56790 2556 56810
rect 2642 56790 2698 56810
rect 2784 56790 2840 56810
rect 2926 56790 2982 56810
rect 3068 56790 3124 56810
rect 2500 56754 2522 56790
rect 2522 56754 2556 56790
rect 2642 56754 2646 56790
rect 2646 56754 2698 56790
rect 2784 56754 2822 56790
rect 2822 56754 2840 56790
rect 2926 56754 2946 56790
rect 2946 56754 2982 56790
rect 3068 56754 3070 56790
rect 3070 56754 3124 56790
rect 3210 56754 3266 56810
rect 3352 56790 3408 56810
rect 3494 56790 3550 56810
rect 3636 56790 3692 56810
rect 3778 56790 3834 56810
rect 3920 56790 3976 56810
rect 3352 56754 3390 56790
rect 3390 56754 3408 56790
rect 3494 56754 3514 56790
rect 3514 56754 3550 56790
rect 3636 56754 3638 56790
rect 3638 56754 3690 56790
rect 3690 56754 3692 56790
rect 3778 56754 3814 56790
rect 3814 56754 3834 56790
rect 3920 56754 3938 56790
rect 3938 56754 3976 56790
rect 4062 56754 4118 56810
rect 4204 56790 4260 56810
rect 4346 56790 4402 56810
rect 4488 56790 4544 56810
rect 4630 56790 4686 56810
rect 4772 56790 4828 56810
rect 4914 56790 4970 56810
rect 4204 56754 4258 56790
rect 4258 56754 4260 56790
rect 4346 56754 4382 56790
rect 4382 56754 4402 56790
rect 4488 56754 4506 56790
rect 4506 56754 4544 56790
rect 4630 56754 4682 56790
rect 4682 56754 4686 56790
rect 4772 56754 4806 56790
rect 4806 56754 4828 56790
rect 4914 56754 4930 56790
rect 4930 56754 4970 56790
rect 5056 56754 5112 56810
rect 5198 56790 5254 56810
rect 5340 56790 5396 56810
rect 5482 56790 5538 56810
rect 5624 56790 5680 56810
rect 5766 56790 5822 56810
rect 5908 56790 5964 56810
rect 5198 56754 5250 56790
rect 5250 56754 5254 56790
rect 5340 56754 5374 56790
rect 5374 56754 5396 56790
rect 5482 56754 5498 56790
rect 5498 56754 5538 56790
rect 5624 56754 5674 56790
rect 5674 56754 5680 56790
rect 5766 56754 5798 56790
rect 5798 56754 5822 56790
rect 5908 56754 5922 56790
rect 5922 56754 5964 56790
rect 6050 56754 6106 56810
rect 6192 56790 6248 56810
rect 6334 56790 6390 56810
rect 6476 56790 6532 56810
rect 6618 56790 6674 56810
rect 6760 56790 6816 56810
rect 6902 56790 6958 56810
rect 6192 56754 6242 56790
rect 6242 56754 6248 56790
rect 6334 56754 6366 56790
rect 6366 56754 6390 56790
rect 6476 56754 6490 56790
rect 6490 56754 6532 56790
rect 6618 56754 6666 56790
rect 6666 56754 6674 56790
rect 6760 56754 6790 56790
rect 6790 56754 6816 56790
rect 6902 56754 6914 56790
rect 6914 56754 6958 56790
rect 7044 56754 7100 56810
rect 7186 56790 7242 56810
rect 7328 56790 7384 56810
rect 7470 56790 7526 56810
rect 7612 56790 7668 56810
rect 7754 56790 7810 56810
rect 7896 56790 7952 56810
rect 7186 56754 7234 56790
rect 7234 56754 7242 56790
rect 7328 56754 7358 56790
rect 7358 56754 7384 56790
rect 7470 56754 7482 56790
rect 7482 56754 7526 56790
rect 7612 56754 7658 56790
rect 7658 56754 7668 56790
rect 7754 56754 7782 56790
rect 7782 56754 7810 56790
rect 7896 56754 7906 56790
rect 7906 56754 7952 56790
rect 8038 56754 8094 56810
rect 8180 56790 8236 56810
rect 8322 56790 8378 56810
rect 8464 56790 8520 56810
rect 8606 56790 8662 56810
rect 8748 56790 8804 56810
rect 8890 56790 8946 56810
rect 8180 56754 8226 56790
rect 8226 56754 8236 56790
rect 8322 56754 8350 56790
rect 8350 56754 8378 56790
rect 8464 56754 8474 56790
rect 8474 56754 8520 56790
rect 8606 56754 8650 56790
rect 8650 56754 8662 56790
rect 8748 56754 8774 56790
rect 8774 56754 8804 56790
rect 8890 56754 8898 56790
rect 8898 56754 8946 56790
rect 9032 56754 9088 56810
rect 9174 56790 9230 56810
rect 9316 56790 9372 56810
rect 9458 56790 9514 56810
rect 9600 56790 9656 56810
rect 9742 56790 9798 56810
rect 9884 56790 9940 56810
rect 9174 56754 9218 56790
rect 9218 56754 9230 56790
rect 9316 56754 9342 56790
rect 9342 56754 9372 56790
rect 9458 56754 9466 56790
rect 9466 56754 9514 56790
rect 9600 56754 9642 56790
rect 9642 56754 9656 56790
rect 9742 56754 9766 56790
rect 9766 56754 9798 56790
rect 9884 56754 9890 56790
rect 9890 56754 9940 56790
rect 10026 56754 10082 56810
rect 10168 56790 10224 56810
rect 10310 56790 10366 56810
rect 10452 56790 10508 56810
rect 10594 56790 10650 56810
rect 10736 56790 10792 56810
rect 10878 56790 10934 56810
rect 10168 56754 10210 56790
rect 10210 56754 10224 56790
rect 10310 56754 10334 56790
rect 10334 56754 10366 56790
rect 10452 56754 10458 56790
rect 10458 56754 10508 56790
rect 10594 56754 10634 56790
rect 10634 56754 10650 56790
rect 10736 56754 10758 56790
rect 10758 56754 10792 56790
rect 10878 56754 10882 56790
rect 10882 56754 10934 56790
rect 11020 56754 11076 56810
rect 11162 56790 11218 56810
rect 11304 56790 11360 56810
rect 11446 56790 11502 56810
rect 11588 56790 11644 56810
rect 11730 56790 11786 56810
rect 11872 56790 11928 56810
rect 11162 56754 11202 56790
rect 11202 56754 11218 56790
rect 11304 56754 11326 56790
rect 11326 56754 11360 56790
rect 11446 56754 11450 56790
rect 11450 56754 11502 56790
rect 11588 56754 11626 56790
rect 11626 56754 11644 56790
rect 11730 56754 11750 56790
rect 11750 56754 11786 56790
rect 11872 56754 11874 56790
rect 11874 56754 11928 56790
rect 12014 56754 12070 56810
rect 12156 56790 12212 56810
rect 12298 56790 12354 56810
rect 12440 56790 12496 56810
rect 12582 56790 12638 56810
rect 12724 56790 12780 56810
rect 12156 56754 12194 56790
rect 12194 56754 12212 56790
rect 12298 56754 12318 56790
rect 12318 56754 12354 56790
rect 12440 56754 12442 56790
rect 12442 56754 12494 56790
rect 12494 56754 12496 56790
rect 12582 56754 12618 56790
rect 12618 56754 12638 56790
rect 12724 56754 12742 56790
rect 12742 56754 12780 56790
rect 12866 56754 12922 56810
rect 13008 56790 13064 56810
rect 13150 56790 13206 56810
rect 13292 56790 13348 56810
rect 13434 56790 13490 56810
rect 13576 56790 13632 56810
rect 13008 56754 13062 56790
rect 13062 56754 13064 56790
rect 13150 56754 13186 56790
rect 13186 56754 13206 56790
rect 13292 56754 13310 56790
rect 13310 56754 13348 56790
rect 13434 56754 13486 56790
rect 13486 56754 13490 56790
rect 13576 56754 13610 56790
rect 13610 56754 13632 56790
rect 2500 56666 2556 56668
rect 2642 56666 2698 56668
rect 2784 56666 2840 56668
rect 2926 56666 2982 56668
rect 3068 56666 3124 56668
rect 2500 56614 2522 56666
rect 2522 56614 2556 56666
rect 2642 56614 2646 56666
rect 2646 56614 2698 56666
rect 2784 56614 2822 56666
rect 2822 56614 2840 56666
rect 2926 56614 2946 56666
rect 2946 56614 2982 56666
rect 3068 56614 3070 56666
rect 3070 56614 3124 56666
rect 2500 56612 2556 56614
rect 2642 56612 2698 56614
rect 2784 56612 2840 56614
rect 2926 56612 2982 56614
rect 3068 56612 3124 56614
rect 3210 56612 3266 56668
rect 3352 56666 3408 56668
rect 3494 56666 3550 56668
rect 3636 56666 3692 56668
rect 3778 56666 3834 56668
rect 3920 56666 3976 56668
rect 3352 56614 3390 56666
rect 3390 56614 3408 56666
rect 3494 56614 3514 56666
rect 3514 56614 3550 56666
rect 3636 56614 3638 56666
rect 3638 56614 3690 56666
rect 3690 56614 3692 56666
rect 3778 56614 3814 56666
rect 3814 56614 3834 56666
rect 3920 56614 3938 56666
rect 3938 56614 3976 56666
rect 3352 56612 3408 56614
rect 3494 56612 3550 56614
rect 3636 56612 3692 56614
rect 3778 56612 3834 56614
rect 3920 56612 3976 56614
rect 4062 56612 4118 56668
rect 4204 56666 4260 56668
rect 4346 56666 4402 56668
rect 4488 56666 4544 56668
rect 4630 56666 4686 56668
rect 4772 56666 4828 56668
rect 4914 56666 4970 56668
rect 4204 56614 4258 56666
rect 4258 56614 4260 56666
rect 4346 56614 4382 56666
rect 4382 56614 4402 56666
rect 4488 56614 4506 56666
rect 4506 56614 4544 56666
rect 4630 56614 4682 56666
rect 4682 56614 4686 56666
rect 4772 56614 4806 56666
rect 4806 56614 4828 56666
rect 4914 56614 4930 56666
rect 4930 56614 4970 56666
rect 4204 56612 4260 56614
rect 4346 56612 4402 56614
rect 4488 56612 4544 56614
rect 4630 56612 4686 56614
rect 4772 56612 4828 56614
rect 4914 56612 4970 56614
rect 5056 56612 5112 56668
rect 5198 56666 5254 56668
rect 5340 56666 5396 56668
rect 5482 56666 5538 56668
rect 5624 56666 5680 56668
rect 5766 56666 5822 56668
rect 5908 56666 5964 56668
rect 5198 56614 5250 56666
rect 5250 56614 5254 56666
rect 5340 56614 5374 56666
rect 5374 56614 5396 56666
rect 5482 56614 5498 56666
rect 5498 56614 5538 56666
rect 5624 56614 5674 56666
rect 5674 56614 5680 56666
rect 5766 56614 5798 56666
rect 5798 56614 5822 56666
rect 5908 56614 5922 56666
rect 5922 56614 5964 56666
rect 5198 56612 5254 56614
rect 5340 56612 5396 56614
rect 5482 56612 5538 56614
rect 5624 56612 5680 56614
rect 5766 56612 5822 56614
rect 5908 56612 5964 56614
rect 6050 56612 6106 56668
rect 6192 56666 6248 56668
rect 6334 56666 6390 56668
rect 6476 56666 6532 56668
rect 6618 56666 6674 56668
rect 6760 56666 6816 56668
rect 6902 56666 6958 56668
rect 6192 56614 6242 56666
rect 6242 56614 6248 56666
rect 6334 56614 6366 56666
rect 6366 56614 6390 56666
rect 6476 56614 6490 56666
rect 6490 56614 6532 56666
rect 6618 56614 6666 56666
rect 6666 56614 6674 56666
rect 6760 56614 6790 56666
rect 6790 56614 6816 56666
rect 6902 56614 6914 56666
rect 6914 56614 6958 56666
rect 6192 56612 6248 56614
rect 6334 56612 6390 56614
rect 6476 56612 6532 56614
rect 6618 56612 6674 56614
rect 6760 56612 6816 56614
rect 6902 56612 6958 56614
rect 7044 56612 7100 56668
rect 7186 56666 7242 56668
rect 7328 56666 7384 56668
rect 7470 56666 7526 56668
rect 7612 56666 7668 56668
rect 7754 56666 7810 56668
rect 7896 56666 7952 56668
rect 7186 56614 7234 56666
rect 7234 56614 7242 56666
rect 7328 56614 7358 56666
rect 7358 56614 7384 56666
rect 7470 56614 7482 56666
rect 7482 56614 7526 56666
rect 7612 56614 7658 56666
rect 7658 56614 7668 56666
rect 7754 56614 7782 56666
rect 7782 56614 7810 56666
rect 7896 56614 7906 56666
rect 7906 56614 7952 56666
rect 7186 56612 7242 56614
rect 7328 56612 7384 56614
rect 7470 56612 7526 56614
rect 7612 56612 7668 56614
rect 7754 56612 7810 56614
rect 7896 56612 7952 56614
rect 8038 56612 8094 56668
rect 8180 56666 8236 56668
rect 8322 56666 8378 56668
rect 8464 56666 8520 56668
rect 8606 56666 8662 56668
rect 8748 56666 8804 56668
rect 8890 56666 8946 56668
rect 8180 56614 8226 56666
rect 8226 56614 8236 56666
rect 8322 56614 8350 56666
rect 8350 56614 8378 56666
rect 8464 56614 8474 56666
rect 8474 56614 8520 56666
rect 8606 56614 8650 56666
rect 8650 56614 8662 56666
rect 8748 56614 8774 56666
rect 8774 56614 8804 56666
rect 8890 56614 8898 56666
rect 8898 56614 8946 56666
rect 8180 56612 8236 56614
rect 8322 56612 8378 56614
rect 8464 56612 8520 56614
rect 8606 56612 8662 56614
rect 8748 56612 8804 56614
rect 8890 56612 8946 56614
rect 9032 56612 9088 56668
rect 9174 56666 9230 56668
rect 9316 56666 9372 56668
rect 9458 56666 9514 56668
rect 9600 56666 9656 56668
rect 9742 56666 9798 56668
rect 9884 56666 9940 56668
rect 9174 56614 9218 56666
rect 9218 56614 9230 56666
rect 9316 56614 9342 56666
rect 9342 56614 9372 56666
rect 9458 56614 9466 56666
rect 9466 56614 9514 56666
rect 9600 56614 9642 56666
rect 9642 56614 9656 56666
rect 9742 56614 9766 56666
rect 9766 56614 9798 56666
rect 9884 56614 9890 56666
rect 9890 56614 9940 56666
rect 9174 56612 9230 56614
rect 9316 56612 9372 56614
rect 9458 56612 9514 56614
rect 9600 56612 9656 56614
rect 9742 56612 9798 56614
rect 9884 56612 9940 56614
rect 10026 56612 10082 56668
rect 10168 56666 10224 56668
rect 10310 56666 10366 56668
rect 10452 56666 10508 56668
rect 10594 56666 10650 56668
rect 10736 56666 10792 56668
rect 10878 56666 10934 56668
rect 10168 56614 10210 56666
rect 10210 56614 10224 56666
rect 10310 56614 10334 56666
rect 10334 56614 10366 56666
rect 10452 56614 10458 56666
rect 10458 56614 10508 56666
rect 10594 56614 10634 56666
rect 10634 56614 10650 56666
rect 10736 56614 10758 56666
rect 10758 56614 10792 56666
rect 10878 56614 10882 56666
rect 10882 56614 10934 56666
rect 10168 56612 10224 56614
rect 10310 56612 10366 56614
rect 10452 56612 10508 56614
rect 10594 56612 10650 56614
rect 10736 56612 10792 56614
rect 10878 56612 10934 56614
rect 11020 56612 11076 56668
rect 11162 56666 11218 56668
rect 11304 56666 11360 56668
rect 11446 56666 11502 56668
rect 11588 56666 11644 56668
rect 11730 56666 11786 56668
rect 11872 56666 11928 56668
rect 11162 56614 11202 56666
rect 11202 56614 11218 56666
rect 11304 56614 11326 56666
rect 11326 56614 11360 56666
rect 11446 56614 11450 56666
rect 11450 56614 11502 56666
rect 11588 56614 11626 56666
rect 11626 56614 11644 56666
rect 11730 56614 11750 56666
rect 11750 56614 11786 56666
rect 11872 56614 11874 56666
rect 11874 56614 11928 56666
rect 11162 56612 11218 56614
rect 11304 56612 11360 56614
rect 11446 56612 11502 56614
rect 11588 56612 11644 56614
rect 11730 56612 11786 56614
rect 11872 56612 11928 56614
rect 12014 56612 12070 56668
rect 12156 56666 12212 56668
rect 12298 56666 12354 56668
rect 12440 56666 12496 56668
rect 12582 56666 12638 56668
rect 12724 56666 12780 56668
rect 12156 56614 12194 56666
rect 12194 56614 12212 56666
rect 12298 56614 12318 56666
rect 12318 56614 12354 56666
rect 12440 56614 12442 56666
rect 12442 56614 12494 56666
rect 12494 56614 12496 56666
rect 12582 56614 12618 56666
rect 12618 56614 12638 56666
rect 12724 56614 12742 56666
rect 12742 56614 12780 56666
rect 12156 56612 12212 56614
rect 12298 56612 12354 56614
rect 12440 56612 12496 56614
rect 12582 56612 12638 56614
rect 12724 56612 12780 56614
rect 12866 56612 12922 56668
rect 13008 56666 13064 56668
rect 13150 56666 13206 56668
rect 13292 56666 13348 56668
rect 13434 56666 13490 56668
rect 13576 56666 13632 56668
rect 13008 56614 13062 56666
rect 13062 56614 13064 56666
rect 13150 56614 13186 56666
rect 13186 56614 13206 56666
rect 13292 56614 13310 56666
rect 13310 56614 13348 56666
rect 13434 56614 13486 56666
rect 13486 56614 13490 56666
rect 13576 56614 13610 56666
rect 13610 56614 13632 56666
rect 13008 56612 13064 56614
rect 13150 56612 13206 56614
rect 13292 56612 13348 56614
rect 13434 56612 13490 56614
rect 13576 56612 13632 56614
rect 2500 56490 2522 56526
rect 2522 56490 2556 56526
rect 2642 56490 2646 56526
rect 2646 56490 2698 56526
rect 2784 56490 2822 56526
rect 2822 56490 2840 56526
rect 2926 56490 2946 56526
rect 2946 56490 2982 56526
rect 3068 56490 3070 56526
rect 3070 56490 3124 56526
rect 2500 56470 2556 56490
rect 2642 56470 2698 56490
rect 2784 56470 2840 56490
rect 2926 56470 2982 56490
rect 3068 56470 3124 56490
rect 3210 56470 3266 56526
rect 3352 56490 3390 56526
rect 3390 56490 3408 56526
rect 3494 56490 3514 56526
rect 3514 56490 3550 56526
rect 3636 56490 3638 56526
rect 3638 56490 3690 56526
rect 3690 56490 3692 56526
rect 3778 56490 3814 56526
rect 3814 56490 3834 56526
rect 3920 56490 3938 56526
rect 3938 56490 3976 56526
rect 3352 56470 3408 56490
rect 3494 56470 3550 56490
rect 3636 56470 3692 56490
rect 3778 56470 3834 56490
rect 3920 56470 3976 56490
rect 4062 56470 4118 56526
rect 4204 56490 4258 56526
rect 4258 56490 4260 56526
rect 4346 56490 4382 56526
rect 4382 56490 4402 56526
rect 4488 56490 4506 56526
rect 4506 56490 4544 56526
rect 4630 56490 4682 56526
rect 4682 56490 4686 56526
rect 4772 56490 4806 56526
rect 4806 56490 4828 56526
rect 4914 56490 4930 56526
rect 4930 56490 4970 56526
rect 4204 56470 4260 56490
rect 4346 56470 4402 56490
rect 4488 56470 4544 56490
rect 4630 56470 4686 56490
rect 4772 56470 4828 56490
rect 4914 56470 4970 56490
rect 5056 56470 5112 56526
rect 5198 56490 5250 56526
rect 5250 56490 5254 56526
rect 5340 56490 5374 56526
rect 5374 56490 5396 56526
rect 5482 56490 5498 56526
rect 5498 56490 5538 56526
rect 5624 56490 5674 56526
rect 5674 56490 5680 56526
rect 5766 56490 5798 56526
rect 5798 56490 5822 56526
rect 5908 56490 5922 56526
rect 5922 56490 5964 56526
rect 5198 56470 5254 56490
rect 5340 56470 5396 56490
rect 5482 56470 5538 56490
rect 5624 56470 5680 56490
rect 5766 56470 5822 56490
rect 5908 56470 5964 56490
rect 6050 56470 6106 56526
rect 6192 56490 6242 56526
rect 6242 56490 6248 56526
rect 6334 56490 6366 56526
rect 6366 56490 6390 56526
rect 6476 56490 6490 56526
rect 6490 56490 6532 56526
rect 6618 56490 6666 56526
rect 6666 56490 6674 56526
rect 6760 56490 6790 56526
rect 6790 56490 6816 56526
rect 6902 56490 6914 56526
rect 6914 56490 6958 56526
rect 6192 56470 6248 56490
rect 6334 56470 6390 56490
rect 6476 56470 6532 56490
rect 6618 56470 6674 56490
rect 6760 56470 6816 56490
rect 6902 56470 6958 56490
rect 7044 56470 7100 56526
rect 7186 56490 7234 56526
rect 7234 56490 7242 56526
rect 7328 56490 7358 56526
rect 7358 56490 7384 56526
rect 7470 56490 7482 56526
rect 7482 56490 7526 56526
rect 7612 56490 7658 56526
rect 7658 56490 7668 56526
rect 7754 56490 7782 56526
rect 7782 56490 7810 56526
rect 7896 56490 7906 56526
rect 7906 56490 7952 56526
rect 7186 56470 7242 56490
rect 7328 56470 7384 56490
rect 7470 56470 7526 56490
rect 7612 56470 7668 56490
rect 7754 56470 7810 56490
rect 7896 56470 7952 56490
rect 8038 56470 8094 56526
rect 8180 56490 8226 56526
rect 8226 56490 8236 56526
rect 8322 56490 8350 56526
rect 8350 56490 8378 56526
rect 8464 56490 8474 56526
rect 8474 56490 8520 56526
rect 8606 56490 8650 56526
rect 8650 56490 8662 56526
rect 8748 56490 8774 56526
rect 8774 56490 8804 56526
rect 8890 56490 8898 56526
rect 8898 56490 8946 56526
rect 8180 56470 8236 56490
rect 8322 56470 8378 56490
rect 8464 56470 8520 56490
rect 8606 56470 8662 56490
rect 8748 56470 8804 56490
rect 8890 56470 8946 56490
rect 9032 56470 9088 56526
rect 9174 56490 9218 56526
rect 9218 56490 9230 56526
rect 9316 56490 9342 56526
rect 9342 56490 9372 56526
rect 9458 56490 9466 56526
rect 9466 56490 9514 56526
rect 9600 56490 9642 56526
rect 9642 56490 9656 56526
rect 9742 56490 9766 56526
rect 9766 56490 9798 56526
rect 9884 56490 9890 56526
rect 9890 56490 9940 56526
rect 9174 56470 9230 56490
rect 9316 56470 9372 56490
rect 9458 56470 9514 56490
rect 9600 56470 9656 56490
rect 9742 56470 9798 56490
rect 9884 56470 9940 56490
rect 10026 56470 10082 56526
rect 10168 56490 10210 56526
rect 10210 56490 10224 56526
rect 10310 56490 10334 56526
rect 10334 56490 10366 56526
rect 10452 56490 10458 56526
rect 10458 56490 10508 56526
rect 10594 56490 10634 56526
rect 10634 56490 10650 56526
rect 10736 56490 10758 56526
rect 10758 56490 10792 56526
rect 10878 56490 10882 56526
rect 10882 56490 10934 56526
rect 10168 56470 10224 56490
rect 10310 56470 10366 56490
rect 10452 56470 10508 56490
rect 10594 56470 10650 56490
rect 10736 56470 10792 56490
rect 10878 56470 10934 56490
rect 11020 56470 11076 56526
rect 11162 56490 11202 56526
rect 11202 56490 11218 56526
rect 11304 56490 11326 56526
rect 11326 56490 11360 56526
rect 11446 56490 11450 56526
rect 11450 56490 11502 56526
rect 11588 56490 11626 56526
rect 11626 56490 11644 56526
rect 11730 56490 11750 56526
rect 11750 56490 11786 56526
rect 11872 56490 11874 56526
rect 11874 56490 11928 56526
rect 11162 56470 11218 56490
rect 11304 56470 11360 56490
rect 11446 56470 11502 56490
rect 11588 56470 11644 56490
rect 11730 56470 11786 56490
rect 11872 56470 11928 56490
rect 12014 56470 12070 56526
rect 12156 56490 12194 56526
rect 12194 56490 12212 56526
rect 12298 56490 12318 56526
rect 12318 56490 12354 56526
rect 12440 56490 12442 56526
rect 12442 56490 12494 56526
rect 12494 56490 12496 56526
rect 12582 56490 12618 56526
rect 12618 56490 12638 56526
rect 12724 56490 12742 56526
rect 12742 56490 12780 56526
rect 12156 56470 12212 56490
rect 12298 56470 12354 56490
rect 12440 56470 12496 56490
rect 12582 56470 12638 56490
rect 12724 56470 12780 56490
rect 12866 56470 12922 56526
rect 13008 56490 13062 56526
rect 13062 56490 13064 56526
rect 13150 56490 13186 56526
rect 13186 56490 13206 56526
rect 13292 56490 13310 56526
rect 13310 56490 13348 56526
rect 13434 56490 13486 56526
rect 13486 56490 13490 56526
rect 13576 56490 13610 56526
rect 13610 56490 13632 56526
rect 13008 56470 13064 56490
rect 13150 56470 13206 56490
rect 13292 56470 13348 56490
rect 13434 56470 13490 56490
rect 13576 56470 13632 56490
rect 2500 56048 2556 56068
rect 2642 56048 2698 56068
rect 2784 56048 2840 56068
rect 2926 56048 2982 56068
rect 3068 56048 3124 56068
rect 2500 56012 2522 56048
rect 2522 56012 2556 56048
rect 2642 56012 2646 56048
rect 2646 56012 2698 56048
rect 2784 56012 2822 56048
rect 2822 56012 2840 56048
rect 2926 56012 2946 56048
rect 2946 56012 2982 56048
rect 3068 56012 3070 56048
rect 3070 56012 3124 56048
rect 3210 56012 3266 56068
rect 3352 56048 3408 56068
rect 3494 56048 3550 56068
rect 3636 56048 3692 56068
rect 3778 56048 3834 56068
rect 3920 56048 3976 56068
rect 3352 56012 3390 56048
rect 3390 56012 3408 56048
rect 3494 56012 3514 56048
rect 3514 56012 3550 56048
rect 3636 56012 3638 56048
rect 3638 56012 3690 56048
rect 3690 56012 3692 56048
rect 3778 56012 3814 56048
rect 3814 56012 3834 56048
rect 3920 56012 3938 56048
rect 3938 56012 3976 56048
rect 4062 56012 4118 56068
rect 4204 56048 4260 56068
rect 4346 56048 4402 56068
rect 4488 56048 4544 56068
rect 4630 56048 4686 56068
rect 4772 56048 4828 56068
rect 4914 56048 4970 56068
rect 4204 56012 4258 56048
rect 4258 56012 4260 56048
rect 4346 56012 4382 56048
rect 4382 56012 4402 56048
rect 4488 56012 4506 56048
rect 4506 56012 4544 56048
rect 4630 56012 4682 56048
rect 4682 56012 4686 56048
rect 4772 56012 4806 56048
rect 4806 56012 4828 56048
rect 4914 56012 4930 56048
rect 4930 56012 4970 56048
rect 5056 56012 5112 56068
rect 5198 56048 5254 56068
rect 5340 56048 5396 56068
rect 5482 56048 5538 56068
rect 5624 56048 5680 56068
rect 5766 56048 5822 56068
rect 5908 56048 5964 56068
rect 5198 56012 5250 56048
rect 5250 56012 5254 56048
rect 5340 56012 5374 56048
rect 5374 56012 5396 56048
rect 5482 56012 5498 56048
rect 5498 56012 5538 56048
rect 5624 56012 5674 56048
rect 5674 56012 5680 56048
rect 5766 56012 5798 56048
rect 5798 56012 5822 56048
rect 5908 56012 5922 56048
rect 5922 56012 5964 56048
rect 6050 56012 6106 56068
rect 6192 56048 6248 56068
rect 6334 56048 6390 56068
rect 6476 56048 6532 56068
rect 6618 56048 6674 56068
rect 6760 56048 6816 56068
rect 6902 56048 6958 56068
rect 6192 56012 6242 56048
rect 6242 56012 6248 56048
rect 6334 56012 6366 56048
rect 6366 56012 6390 56048
rect 6476 56012 6490 56048
rect 6490 56012 6532 56048
rect 6618 56012 6666 56048
rect 6666 56012 6674 56048
rect 6760 56012 6790 56048
rect 6790 56012 6816 56048
rect 6902 56012 6914 56048
rect 6914 56012 6958 56048
rect 7044 56012 7100 56068
rect 7186 56048 7242 56068
rect 7328 56048 7384 56068
rect 7470 56048 7526 56068
rect 7612 56048 7668 56068
rect 7754 56048 7810 56068
rect 7896 56048 7952 56068
rect 7186 56012 7234 56048
rect 7234 56012 7242 56048
rect 7328 56012 7358 56048
rect 7358 56012 7384 56048
rect 7470 56012 7482 56048
rect 7482 56012 7526 56048
rect 7612 56012 7658 56048
rect 7658 56012 7668 56048
rect 7754 56012 7782 56048
rect 7782 56012 7810 56048
rect 7896 56012 7906 56048
rect 7906 56012 7952 56048
rect 8038 56012 8094 56068
rect 8180 56048 8236 56068
rect 8322 56048 8378 56068
rect 8464 56048 8520 56068
rect 8606 56048 8662 56068
rect 8748 56048 8804 56068
rect 8890 56048 8946 56068
rect 8180 56012 8226 56048
rect 8226 56012 8236 56048
rect 8322 56012 8350 56048
rect 8350 56012 8378 56048
rect 8464 56012 8474 56048
rect 8474 56012 8520 56048
rect 8606 56012 8650 56048
rect 8650 56012 8662 56048
rect 8748 56012 8774 56048
rect 8774 56012 8804 56048
rect 8890 56012 8898 56048
rect 8898 56012 8946 56048
rect 9032 56012 9088 56068
rect 9174 56048 9230 56068
rect 9316 56048 9372 56068
rect 9458 56048 9514 56068
rect 9600 56048 9656 56068
rect 9742 56048 9798 56068
rect 9884 56048 9940 56068
rect 9174 56012 9218 56048
rect 9218 56012 9230 56048
rect 9316 56012 9342 56048
rect 9342 56012 9372 56048
rect 9458 56012 9466 56048
rect 9466 56012 9514 56048
rect 9600 56012 9642 56048
rect 9642 56012 9656 56048
rect 9742 56012 9766 56048
rect 9766 56012 9798 56048
rect 9884 56012 9890 56048
rect 9890 56012 9940 56048
rect 10026 56012 10082 56068
rect 10168 56048 10224 56068
rect 10310 56048 10366 56068
rect 10452 56048 10508 56068
rect 10594 56048 10650 56068
rect 10736 56048 10792 56068
rect 10878 56048 10934 56068
rect 10168 56012 10210 56048
rect 10210 56012 10224 56048
rect 10310 56012 10334 56048
rect 10334 56012 10366 56048
rect 10452 56012 10458 56048
rect 10458 56012 10508 56048
rect 10594 56012 10634 56048
rect 10634 56012 10650 56048
rect 10736 56012 10758 56048
rect 10758 56012 10792 56048
rect 10878 56012 10882 56048
rect 10882 56012 10934 56048
rect 11020 56012 11076 56068
rect 11162 56048 11218 56068
rect 11304 56048 11360 56068
rect 11446 56048 11502 56068
rect 11588 56048 11644 56068
rect 11730 56048 11786 56068
rect 11872 56048 11928 56068
rect 11162 56012 11202 56048
rect 11202 56012 11218 56048
rect 11304 56012 11326 56048
rect 11326 56012 11360 56048
rect 11446 56012 11450 56048
rect 11450 56012 11502 56048
rect 11588 56012 11626 56048
rect 11626 56012 11644 56048
rect 11730 56012 11750 56048
rect 11750 56012 11786 56048
rect 11872 56012 11874 56048
rect 11874 56012 11928 56048
rect 12014 56012 12070 56068
rect 12156 56048 12212 56068
rect 12298 56048 12354 56068
rect 12440 56048 12496 56068
rect 12582 56048 12638 56068
rect 12724 56048 12780 56068
rect 12156 56012 12194 56048
rect 12194 56012 12212 56048
rect 12298 56012 12318 56048
rect 12318 56012 12354 56048
rect 12440 56012 12442 56048
rect 12442 56012 12494 56048
rect 12494 56012 12496 56048
rect 12582 56012 12618 56048
rect 12618 56012 12638 56048
rect 12724 56012 12742 56048
rect 12742 56012 12780 56048
rect 12866 56012 12922 56068
rect 13008 56048 13064 56068
rect 13150 56048 13206 56068
rect 13292 56048 13348 56068
rect 13434 56048 13490 56068
rect 13576 56048 13632 56068
rect 13008 56012 13062 56048
rect 13062 56012 13064 56048
rect 13150 56012 13186 56048
rect 13186 56012 13206 56048
rect 13292 56012 13310 56048
rect 13310 56012 13348 56048
rect 13434 56012 13486 56048
rect 13486 56012 13490 56048
rect 13576 56012 13610 56048
rect 13610 56012 13632 56048
rect 2500 55924 2556 55926
rect 2642 55924 2698 55926
rect 2784 55924 2840 55926
rect 2926 55924 2982 55926
rect 3068 55924 3124 55926
rect 2500 55872 2522 55924
rect 2522 55872 2556 55924
rect 2642 55872 2646 55924
rect 2646 55872 2698 55924
rect 2784 55872 2822 55924
rect 2822 55872 2840 55924
rect 2926 55872 2946 55924
rect 2946 55872 2982 55924
rect 3068 55872 3070 55924
rect 3070 55872 3124 55924
rect 2500 55870 2556 55872
rect 2642 55870 2698 55872
rect 2784 55870 2840 55872
rect 2926 55870 2982 55872
rect 3068 55870 3124 55872
rect 3210 55870 3266 55926
rect 3352 55924 3408 55926
rect 3494 55924 3550 55926
rect 3636 55924 3692 55926
rect 3778 55924 3834 55926
rect 3920 55924 3976 55926
rect 3352 55872 3390 55924
rect 3390 55872 3408 55924
rect 3494 55872 3514 55924
rect 3514 55872 3550 55924
rect 3636 55872 3638 55924
rect 3638 55872 3690 55924
rect 3690 55872 3692 55924
rect 3778 55872 3814 55924
rect 3814 55872 3834 55924
rect 3920 55872 3938 55924
rect 3938 55872 3976 55924
rect 3352 55870 3408 55872
rect 3494 55870 3550 55872
rect 3636 55870 3692 55872
rect 3778 55870 3834 55872
rect 3920 55870 3976 55872
rect 4062 55870 4118 55926
rect 4204 55924 4260 55926
rect 4346 55924 4402 55926
rect 4488 55924 4544 55926
rect 4630 55924 4686 55926
rect 4772 55924 4828 55926
rect 4914 55924 4970 55926
rect 4204 55872 4258 55924
rect 4258 55872 4260 55924
rect 4346 55872 4382 55924
rect 4382 55872 4402 55924
rect 4488 55872 4506 55924
rect 4506 55872 4544 55924
rect 4630 55872 4682 55924
rect 4682 55872 4686 55924
rect 4772 55872 4806 55924
rect 4806 55872 4828 55924
rect 4914 55872 4930 55924
rect 4930 55872 4970 55924
rect 4204 55870 4260 55872
rect 4346 55870 4402 55872
rect 4488 55870 4544 55872
rect 4630 55870 4686 55872
rect 4772 55870 4828 55872
rect 4914 55870 4970 55872
rect 5056 55870 5112 55926
rect 5198 55924 5254 55926
rect 5340 55924 5396 55926
rect 5482 55924 5538 55926
rect 5624 55924 5680 55926
rect 5766 55924 5822 55926
rect 5908 55924 5964 55926
rect 5198 55872 5250 55924
rect 5250 55872 5254 55924
rect 5340 55872 5374 55924
rect 5374 55872 5396 55924
rect 5482 55872 5498 55924
rect 5498 55872 5538 55924
rect 5624 55872 5674 55924
rect 5674 55872 5680 55924
rect 5766 55872 5798 55924
rect 5798 55872 5822 55924
rect 5908 55872 5922 55924
rect 5922 55872 5964 55924
rect 5198 55870 5254 55872
rect 5340 55870 5396 55872
rect 5482 55870 5538 55872
rect 5624 55870 5680 55872
rect 5766 55870 5822 55872
rect 5908 55870 5964 55872
rect 6050 55870 6106 55926
rect 6192 55924 6248 55926
rect 6334 55924 6390 55926
rect 6476 55924 6532 55926
rect 6618 55924 6674 55926
rect 6760 55924 6816 55926
rect 6902 55924 6958 55926
rect 6192 55872 6242 55924
rect 6242 55872 6248 55924
rect 6334 55872 6366 55924
rect 6366 55872 6390 55924
rect 6476 55872 6490 55924
rect 6490 55872 6532 55924
rect 6618 55872 6666 55924
rect 6666 55872 6674 55924
rect 6760 55872 6790 55924
rect 6790 55872 6816 55924
rect 6902 55872 6914 55924
rect 6914 55872 6958 55924
rect 6192 55870 6248 55872
rect 6334 55870 6390 55872
rect 6476 55870 6532 55872
rect 6618 55870 6674 55872
rect 6760 55870 6816 55872
rect 6902 55870 6958 55872
rect 7044 55870 7100 55926
rect 7186 55924 7242 55926
rect 7328 55924 7384 55926
rect 7470 55924 7526 55926
rect 7612 55924 7668 55926
rect 7754 55924 7810 55926
rect 7896 55924 7952 55926
rect 7186 55872 7234 55924
rect 7234 55872 7242 55924
rect 7328 55872 7358 55924
rect 7358 55872 7384 55924
rect 7470 55872 7482 55924
rect 7482 55872 7526 55924
rect 7612 55872 7658 55924
rect 7658 55872 7668 55924
rect 7754 55872 7782 55924
rect 7782 55872 7810 55924
rect 7896 55872 7906 55924
rect 7906 55872 7952 55924
rect 7186 55870 7242 55872
rect 7328 55870 7384 55872
rect 7470 55870 7526 55872
rect 7612 55870 7668 55872
rect 7754 55870 7810 55872
rect 7896 55870 7952 55872
rect 8038 55870 8094 55926
rect 8180 55924 8236 55926
rect 8322 55924 8378 55926
rect 8464 55924 8520 55926
rect 8606 55924 8662 55926
rect 8748 55924 8804 55926
rect 8890 55924 8946 55926
rect 8180 55872 8226 55924
rect 8226 55872 8236 55924
rect 8322 55872 8350 55924
rect 8350 55872 8378 55924
rect 8464 55872 8474 55924
rect 8474 55872 8520 55924
rect 8606 55872 8650 55924
rect 8650 55872 8662 55924
rect 8748 55872 8774 55924
rect 8774 55872 8804 55924
rect 8890 55872 8898 55924
rect 8898 55872 8946 55924
rect 8180 55870 8236 55872
rect 8322 55870 8378 55872
rect 8464 55870 8520 55872
rect 8606 55870 8662 55872
rect 8748 55870 8804 55872
rect 8890 55870 8946 55872
rect 9032 55870 9088 55926
rect 9174 55924 9230 55926
rect 9316 55924 9372 55926
rect 9458 55924 9514 55926
rect 9600 55924 9656 55926
rect 9742 55924 9798 55926
rect 9884 55924 9940 55926
rect 9174 55872 9218 55924
rect 9218 55872 9230 55924
rect 9316 55872 9342 55924
rect 9342 55872 9372 55924
rect 9458 55872 9466 55924
rect 9466 55872 9514 55924
rect 9600 55872 9642 55924
rect 9642 55872 9656 55924
rect 9742 55872 9766 55924
rect 9766 55872 9798 55924
rect 9884 55872 9890 55924
rect 9890 55872 9940 55924
rect 9174 55870 9230 55872
rect 9316 55870 9372 55872
rect 9458 55870 9514 55872
rect 9600 55870 9656 55872
rect 9742 55870 9798 55872
rect 9884 55870 9940 55872
rect 10026 55870 10082 55926
rect 10168 55924 10224 55926
rect 10310 55924 10366 55926
rect 10452 55924 10508 55926
rect 10594 55924 10650 55926
rect 10736 55924 10792 55926
rect 10878 55924 10934 55926
rect 10168 55872 10210 55924
rect 10210 55872 10224 55924
rect 10310 55872 10334 55924
rect 10334 55872 10366 55924
rect 10452 55872 10458 55924
rect 10458 55872 10508 55924
rect 10594 55872 10634 55924
rect 10634 55872 10650 55924
rect 10736 55872 10758 55924
rect 10758 55872 10792 55924
rect 10878 55872 10882 55924
rect 10882 55872 10934 55924
rect 10168 55870 10224 55872
rect 10310 55870 10366 55872
rect 10452 55870 10508 55872
rect 10594 55870 10650 55872
rect 10736 55870 10792 55872
rect 10878 55870 10934 55872
rect 11020 55870 11076 55926
rect 11162 55924 11218 55926
rect 11304 55924 11360 55926
rect 11446 55924 11502 55926
rect 11588 55924 11644 55926
rect 11730 55924 11786 55926
rect 11872 55924 11928 55926
rect 11162 55872 11202 55924
rect 11202 55872 11218 55924
rect 11304 55872 11326 55924
rect 11326 55872 11360 55924
rect 11446 55872 11450 55924
rect 11450 55872 11502 55924
rect 11588 55872 11626 55924
rect 11626 55872 11644 55924
rect 11730 55872 11750 55924
rect 11750 55872 11786 55924
rect 11872 55872 11874 55924
rect 11874 55872 11928 55924
rect 11162 55870 11218 55872
rect 11304 55870 11360 55872
rect 11446 55870 11502 55872
rect 11588 55870 11644 55872
rect 11730 55870 11786 55872
rect 11872 55870 11928 55872
rect 12014 55870 12070 55926
rect 12156 55924 12212 55926
rect 12298 55924 12354 55926
rect 12440 55924 12496 55926
rect 12582 55924 12638 55926
rect 12724 55924 12780 55926
rect 12156 55872 12194 55924
rect 12194 55872 12212 55924
rect 12298 55872 12318 55924
rect 12318 55872 12354 55924
rect 12440 55872 12442 55924
rect 12442 55872 12494 55924
rect 12494 55872 12496 55924
rect 12582 55872 12618 55924
rect 12618 55872 12638 55924
rect 12724 55872 12742 55924
rect 12742 55872 12780 55924
rect 12156 55870 12212 55872
rect 12298 55870 12354 55872
rect 12440 55870 12496 55872
rect 12582 55870 12638 55872
rect 12724 55870 12780 55872
rect 12866 55870 12922 55926
rect 13008 55924 13064 55926
rect 13150 55924 13206 55926
rect 13292 55924 13348 55926
rect 13434 55924 13490 55926
rect 13576 55924 13632 55926
rect 13008 55872 13062 55924
rect 13062 55872 13064 55924
rect 13150 55872 13186 55924
rect 13186 55872 13206 55924
rect 13292 55872 13310 55924
rect 13310 55872 13348 55924
rect 13434 55872 13486 55924
rect 13486 55872 13490 55924
rect 13576 55872 13610 55924
rect 13610 55872 13632 55924
rect 13008 55870 13064 55872
rect 13150 55870 13206 55872
rect 13292 55870 13348 55872
rect 13434 55870 13490 55872
rect 13576 55870 13632 55872
rect 2500 55748 2522 55784
rect 2522 55748 2556 55784
rect 2642 55748 2646 55784
rect 2646 55748 2698 55784
rect 2784 55748 2822 55784
rect 2822 55748 2840 55784
rect 2926 55748 2946 55784
rect 2946 55748 2982 55784
rect 3068 55748 3070 55784
rect 3070 55748 3124 55784
rect 2500 55728 2556 55748
rect 2642 55728 2698 55748
rect 2784 55728 2840 55748
rect 2926 55728 2982 55748
rect 3068 55728 3124 55748
rect 3210 55728 3266 55784
rect 3352 55748 3390 55784
rect 3390 55748 3408 55784
rect 3494 55748 3514 55784
rect 3514 55748 3550 55784
rect 3636 55748 3638 55784
rect 3638 55748 3690 55784
rect 3690 55748 3692 55784
rect 3778 55748 3814 55784
rect 3814 55748 3834 55784
rect 3920 55748 3938 55784
rect 3938 55748 3976 55784
rect 3352 55728 3408 55748
rect 3494 55728 3550 55748
rect 3636 55728 3692 55748
rect 3778 55728 3834 55748
rect 3920 55728 3976 55748
rect 4062 55728 4118 55784
rect 4204 55748 4258 55784
rect 4258 55748 4260 55784
rect 4346 55748 4382 55784
rect 4382 55748 4402 55784
rect 4488 55748 4506 55784
rect 4506 55748 4544 55784
rect 4630 55748 4682 55784
rect 4682 55748 4686 55784
rect 4772 55748 4806 55784
rect 4806 55748 4828 55784
rect 4914 55748 4930 55784
rect 4930 55748 4970 55784
rect 4204 55728 4260 55748
rect 4346 55728 4402 55748
rect 4488 55728 4544 55748
rect 4630 55728 4686 55748
rect 4772 55728 4828 55748
rect 4914 55728 4970 55748
rect 5056 55728 5112 55784
rect 5198 55748 5250 55784
rect 5250 55748 5254 55784
rect 5340 55748 5374 55784
rect 5374 55748 5396 55784
rect 5482 55748 5498 55784
rect 5498 55748 5538 55784
rect 5624 55748 5674 55784
rect 5674 55748 5680 55784
rect 5766 55748 5798 55784
rect 5798 55748 5822 55784
rect 5908 55748 5922 55784
rect 5922 55748 5964 55784
rect 5198 55728 5254 55748
rect 5340 55728 5396 55748
rect 5482 55728 5538 55748
rect 5624 55728 5680 55748
rect 5766 55728 5822 55748
rect 5908 55728 5964 55748
rect 6050 55728 6106 55784
rect 6192 55748 6242 55784
rect 6242 55748 6248 55784
rect 6334 55748 6366 55784
rect 6366 55748 6390 55784
rect 6476 55748 6490 55784
rect 6490 55748 6532 55784
rect 6618 55748 6666 55784
rect 6666 55748 6674 55784
rect 6760 55748 6790 55784
rect 6790 55748 6816 55784
rect 6902 55748 6914 55784
rect 6914 55748 6958 55784
rect 6192 55728 6248 55748
rect 6334 55728 6390 55748
rect 6476 55728 6532 55748
rect 6618 55728 6674 55748
rect 6760 55728 6816 55748
rect 6902 55728 6958 55748
rect 7044 55728 7100 55784
rect 7186 55748 7234 55784
rect 7234 55748 7242 55784
rect 7328 55748 7358 55784
rect 7358 55748 7384 55784
rect 7470 55748 7482 55784
rect 7482 55748 7526 55784
rect 7612 55748 7658 55784
rect 7658 55748 7668 55784
rect 7754 55748 7782 55784
rect 7782 55748 7810 55784
rect 7896 55748 7906 55784
rect 7906 55748 7952 55784
rect 7186 55728 7242 55748
rect 7328 55728 7384 55748
rect 7470 55728 7526 55748
rect 7612 55728 7668 55748
rect 7754 55728 7810 55748
rect 7896 55728 7952 55748
rect 8038 55728 8094 55784
rect 8180 55748 8226 55784
rect 8226 55748 8236 55784
rect 8322 55748 8350 55784
rect 8350 55748 8378 55784
rect 8464 55748 8474 55784
rect 8474 55748 8520 55784
rect 8606 55748 8650 55784
rect 8650 55748 8662 55784
rect 8748 55748 8774 55784
rect 8774 55748 8804 55784
rect 8890 55748 8898 55784
rect 8898 55748 8946 55784
rect 8180 55728 8236 55748
rect 8322 55728 8378 55748
rect 8464 55728 8520 55748
rect 8606 55728 8662 55748
rect 8748 55728 8804 55748
rect 8890 55728 8946 55748
rect 9032 55728 9088 55784
rect 9174 55748 9218 55784
rect 9218 55748 9230 55784
rect 9316 55748 9342 55784
rect 9342 55748 9372 55784
rect 9458 55748 9466 55784
rect 9466 55748 9514 55784
rect 9600 55748 9642 55784
rect 9642 55748 9656 55784
rect 9742 55748 9766 55784
rect 9766 55748 9798 55784
rect 9884 55748 9890 55784
rect 9890 55748 9940 55784
rect 9174 55728 9230 55748
rect 9316 55728 9372 55748
rect 9458 55728 9514 55748
rect 9600 55728 9656 55748
rect 9742 55728 9798 55748
rect 9884 55728 9940 55748
rect 10026 55728 10082 55784
rect 10168 55748 10210 55784
rect 10210 55748 10224 55784
rect 10310 55748 10334 55784
rect 10334 55748 10366 55784
rect 10452 55748 10458 55784
rect 10458 55748 10508 55784
rect 10594 55748 10634 55784
rect 10634 55748 10650 55784
rect 10736 55748 10758 55784
rect 10758 55748 10792 55784
rect 10878 55748 10882 55784
rect 10882 55748 10934 55784
rect 10168 55728 10224 55748
rect 10310 55728 10366 55748
rect 10452 55728 10508 55748
rect 10594 55728 10650 55748
rect 10736 55728 10792 55748
rect 10878 55728 10934 55748
rect 11020 55728 11076 55784
rect 11162 55748 11202 55784
rect 11202 55748 11218 55784
rect 11304 55748 11326 55784
rect 11326 55748 11360 55784
rect 11446 55748 11450 55784
rect 11450 55748 11502 55784
rect 11588 55748 11626 55784
rect 11626 55748 11644 55784
rect 11730 55748 11750 55784
rect 11750 55748 11786 55784
rect 11872 55748 11874 55784
rect 11874 55748 11928 55784
rect 11162 55728 11218 55748
rect 11304 55728 11360 55748
rect 11446 55728 11502 55748
rect 11588 55728 11644 55748
rect 11730 55728 11786 55748
rect 11872 55728 11928 55748
rect 12014 55728 12070 55784
rect 12156 55748 12194 55784
rect 12194 55748 12212 55784
rect 12298 55748 12318 55784
rect 12318 55748 12354 55784
rect 12440 55748 12442 55784
rect 12442 55748 12494 55784
rect 12494 55748 12496 55784
rect 12582 55748 12618 55784
rect 12618 55748 12638 55784
rect 12724 55748 12742 55784
rect 12742 55748 12780 55784
rect 12156 55728 12212 55748
rect 12298 55728 12354 55748
rect 12440 55728 12496 55748
rect 12582 55728 12638 55748
rect 12724 55728 12780 55748
rect 12866 55728 12922 55784
rect 13008 55748 13062 55784
rect 13062 55748 13064 55784
rect 13150 55748 13186 55784
rect 13186 55748 13206 55784
rect 13292 55748 13310 55784
rect 13310 55748 13348 55784
rect 13434 55748 13486 55784
rect 13486 55748 13490 55784
rect 13576 55748 13610 55784
rect 13610 55748 13632 55784
rect 13008 55728 13064 55748
rect 13150 55728 13206 55748
rect 13292 55728 13348 55748
rect 13434 55728 13490 55748
rect 13576 55728 13632 55748
rect 4768 55341 4770 55397
rect 4770 55341 4822 55397
rect 4822 55341 4824 55397
rect 4768 55199 4770 55255
rect 4770 55199 4822 55255
rect 4822 55199 4824 55255
rect 4768 55057 4770 55113
rect 4770 55057 4822 55113
rect 4822 55057 4824 55113
rect 4768 54915 4770 54971
rect 4770 54915 4822 54971
rect 4822 54915 4824 54971
rect 4768 54773 4770 54829
rect 4770 54773 4822 54829
rect 4822 54773 4824 54829
rect 4768 54631 4770 54687
rect 4770 54631 4822 54687
rect 4822 54631 4824 54687
rect 4948 55341 4950 55397
rect 4950 55341 5002 55397
rect 5002 55341 5004 55397
rect 4948 55199 4950 55255
rect 4950 55199 5002 55255
rect 5002 55199 5004 55255
rect 4948 55057 4950 55113
rect 4950 55057 5002 55113
rect 5002 55057 5004 55113
rect 4948 54915 4950 54971
rect 4950 54915 5002 54971
rect 5002 54915 5004 54971
rect 4948 54773 4950 54829
rect 4950 54773 5002 54829
rect 5002 54773 5004 54829
rect 4948 54631 4950 54687
rect 4950 54631 5002 54687
rect 5002 54631 5004 54687
rect 5436 55341 5438 55397
rect 5438 55341 5490 55397
rect 5490 55341 5492 55397
rect 5436 55199 5438 55255
rect 5438 55199 5490 55255
rect 5490 55199 5492 55255
rect 5436 55057 5438 55113
rect 5438 55057 5490 55113
rect 5490 55057 5492 55113
rect 5436 54915 5438 54971
rect 5438 54915 5490 54971
rect 5490 54915 5492 54971
rect 5436 54773 5438 54829
rect 5438 54773 5490 54829
rect 5490 54773 5492 54829
rect 5436 54631 5438 54687
rect 5438 54631 5490 54687
rect 5490 54631 5492 54687
rect 5924 55341 5926 55397
rect 5926 55341 5978 55397
rect 5978 55341 5980 55397
rect 5924 55199 5926 55255
rect 5926 55199 5978 55255
rect 5978 55199 5980 55255
rect 5924 55057 5926 55113
rect 5926 55057 5978 55113
rect 5978 55057 5980 55113
rect 5924 54915 5926 54971
rect 5926 54915 5978 54971
rect 5978 54915 5980 54971
rect 5924 54773 5926 54829
rect 5926 54773 5978 54829
rect 5978 54773 5980 54829
rect 5924 54631 5926 54687
rect 5926 54631 5978 54687
rect 5978 54631 5980 54687
rect 6106 55359 6162 55371
rect 6106 55315 6108 55359
rect 6108 55315 6160 55359
rect 6160 55315 6162 55359
rect 6106 55173 6108 55229
rect 6108 55173 6160 55229
rect 6160 55173 6162 55229
rect 6106 55031 6108 55087
rect 6108 55031 6160 55087
rect 6160 55031 6162 55087
rect 6106 54889 6108 54945
rect 6108 54889 6160 54945
rect 6160 54889 6162 54945
rect 6106 54747 6108 54803
rect 6108 54747 6160 54803
rect 6160 54747 6162 54803
rect 6106 54605 6108 54661
rect 6108 54605 6160 54661
rect 6160 54605 6162 54661
rect 6288 55341 6290 55397
rect 6290 55341 6342 55397
rect 6342 55341 6344 55397
rect 6288 55199 6290 55255
rect 6290 55199 6342 55255
rect 6342 55199 6344 55255
rect 6288 55057 6290 55113
rect 6290 55057 6342 55113
rect 6342 55057 6344 55113
rect 6288 54915 6290 54971
rect 6290 54915 6342 54971
rect 6342 54915 6344 54971
rect 6288 54773 6290 54829
rect 6290 54773 6342 54829
rect 6342 54773 6344 54829
rect 6288 54631 6290 54687
rect 6290 54631 6342 54687
rect 6342 54631 6344 54687
rect 6776 55341 6778 55397
rect 6778 55341 6830 55397
rect 6830 55341 6832 55397
rect 6776 55199 6778 55255
rect 6778 55199 6830 55255
rect 6830 55199 6832 55255
rect 6776 55057 6778 55113
rect 6778 55057 6830 55113
rect 6830 55057 6832 55113
rect 6776 54915 6778 54971
rect 6778 54915 6830 54971
rect 6830 54915 6832 54971
rect 6776 54773 6778 54829
rect 6778 54773 6830 54829
rect 6830 54773 6832 54829
rect 6776 54631 6778 54687
rect 6778 54631 6830 54687
rect 6830 54631 6832 54687
rect 7264 55341 7266 55397
rect 7266 55341 7318 55397
rect 7318 55341 7320 55397
rect 7264 55199 7266 55255
rect 7266 55199 7318 55255
rect 7318 55199 7320 55255
rect 7264 55057 7266 55113
rect 7266 55057 7318 55113
rect 7318 55057 7320 55113
rect 7264 54915 7266 54971
rect 7266 54915 7318 54971
rect 7318 54915 7320 54971
rect 7264 54773 7266 54829
rect 7266 54773 7318 54829
rect 7318 54773 7320 54829
rect 7264 54631 7266 54687
rect 7266 54631 7318 54687
rect 7318 54631 7320 54687
rect 7444 55341 7446 55397
rect 7446 55341 7498 55397
rect 7498 55341 7500 55397
rect 7444 55199 7446 55255
rect 7446 55199 7498 55255
rect 7498 55199 7500 55255
rect 7444 55057 7446 55113
rect 7446 55057 7498 55113
rect 7498 55057 7500 55113
rect 7444 54915 7446 54971
rect 7446 54915 7498 54971
rect 7498 54915 7500 54971
rect 7444 54773 7446 54829
rect 7446 54773 7498 54829
rect 7498 54773 7500 54829
rect 7444 54631 7446 54687
rect 7446 54631 7498 54687
rect 7498 54631 7500 54687
rect 6106 54475 6108 54519
rect 6108 54475 6160 54519
rect 6160 54475 6162 54519
rect 6106 54463 6162 54475
rect 10012 55341 10014 55397
rect 10014 55341 10066 55397
rect 10066 55341 10068 55397
rect 10012 55199 10014 55255
rect 10014 55199 10066 55255
rect 10066 55199 10068 55255
rect 10012 55057 10014 55113
rect 10014 55057 10066 55113
rect 10066 55057 10068 55113
rect 10012 54915 10014 54971
rect 10014 54915 10066 54971
rect 10066 54915 10068 54971
rect 10012 54773 10014 54829
rect 10014 54773 10066 54829
rect 10066 54773 10068 54829
rect 10012 54631 10014 54687
rect 10014 54631 10066 54687
rect 10066 54631 10068 54687
rect 10192 55341 10194 55397
rect 10194 55341 10246 55397
rect 10246 55341 10248 55397
rect 10192 55199 10194 55255
rect 10194 55199 10246 55255
rect 10246 55199 10248 55255
rect 10192 55057 10194 55113
rect 10194 55057 10246 55113
rect 10246 55057 10248 55113
rect 10192 54915 10194 54971
rect 10194 54915 10246 54971
rect 10246 54915 10248 54971
rect 10192 54773 10194 54829
rect 10194 54773 10246 54829
rect 10246 54773 10248 54829
rect 10192 54631 10194 54687
rect 10194 54631 10246 54687
rect 10246 54631 10248 54687
rect 10680 55341 10682 55397
rect 10682 55341 10734 55397
rect 10734 55341 10736 55397
rect 10680 55199 10682 55255
rect 10682 55199 10734 55255
rect 10734 55199 10736 55255
rect 10680 55057 10682 55113
rect 10682 55057 10734 55113
rect 10734 55057 10736 55113
rect 10680 54915 10682 54971
rect 10682 54915 10734 54971
rect 10734 54915 10736 54971
rect 10680 54773 10682 54829
rect 10682 54773 10734 54829
rect 10734 54773 10736 54829
rect 10680 54631 10682 54687
rect 10682 54631 10734 54687
rect 10734 54631 10736 54687
rect 11168 55341 11170 55397
rect 11170 55341 11222 55397
rect 11222 55341 11224 55397
rect 11168 55199 11170 55255
rect 11170 55199 11222 55255
rect 11222 55199 11224 55255
rect 11168 55057 11170 55113
rect 11170 55057 11222 55113
rect 11222 55057 11224 55113
rect 11168 54915 11170 54971
rect 11170 54915 11222 54971
rect 11222 54915 11224 54971
rect 11168 54773 11170 54829
rect 11170 54773 11222 54829
rect 11222 54773 11224 54829
rect 11168 54631 11170 54687
rect 11170 54631 11222 54687
rect 11222 54631 11224 54687
rect 11350 55359 11406 55371
rect 11350 55315 11352 55359
rect 11352 55315 11404 55359
rect 11404 55315 11406 55359
rect 11350 55173 11352 55229
rect 11352 55173 11404 55229
rect 11404 55173 11406 55229
rect 11350 55031 11352 55087
rect 11352 55031 11404 55087
rect 11404 55031 11406 55087
rect 11350 54889 11352 54945
rect 11352 54889 11404 54945
rect 11404 54889 11406 54945
rect 11350 54747 11352 54803
rect 11352 54747 11404 54803
rect 11404 54747 11406 54803
rect 11350 54605 11352 54661
rect 11352 54605 11404 54661
rect 11404 54605 11406 54661
rect 11532 55341 11534 55397
rect 11534 55341 11586 55397
rect 11586 55341 11588 55397
rect 11532 55199 11534 55255
rect 11534 55199 11586 55255
rect 11586 55199 11588 55255
rect 11532 55057 11534 55113
rect 11534 55057 11586 55113
rect 11586 55057 11588 55113
rect 11532 54915 11534 54971
rect 11534 54915 11586 54971
rect 11586 54915 11588 54971
rect 11532 54773 11534 54829
rect 11534 54773 11586 54829
rect 11586 54773 11588 54829
rect 11532 54631 11534 54687
rect 11534 54631 11586 54687
rect 11586 54631 11588 54687
rect 12020 55341 12022 55397
rect 12022 55341 12074 55397
rect 12074 55341 12076 55397
rect 12020 55199 12022 55255
rect 12022 55199 12074 55255
rect 12074 55199 12076 55255
rect 12020 55057 12022 55113
rect 12022 55057 12074 55113
rect 12074 55057 12076 55113
rect 12020 54915 12022 54971
rect 12022 54915 12074 54971
rect 12074 54915 12076 54971
rect 12020 54773 12022 54829
rect 12022 54773 12074 54829
rect 12074 54773 12076 54829
rect 12020 54631 12022 54687
rect 12022 54631 12074 54687
rect 12074 54631 12076 54687
rect 12508 55341 12510 55397
rect 12510 55341 12562 55397
rect 12562 55341 12564 55397
rect 12508 55199 12510 55255
rect 12510 55199 12562 55255
rect 12562 55199 12564 55255
rect 12508 55057 12510 55113
rect 12510 55057 12562 55113
rect 12562 55057 12564 55113
rect 12508 54915 12510 54971
rect 12510 54915 12562 54971
rect 12562 54915 12564 54971
rect 12508 54773 12510 54829
rect 12510 54773 12562 54829
rect 12562 54773 12564 54829
rect 12508 54631 12510 54687
rect 12510 54631 12562 54687
rect 12562 54631 12564 54687
rect 12688 55341 12690 55397
rect 12690 55341 12742 55397
rect 12742 55341 12744 55397
rect 12688 55199 12690 55255
rect 12690 55199 12742 55255
rect 12742 55199 12744 55255
rect 12688 55057 12690 55113
rect 12690 55057 12742 55113
rect 12742 55057 12744 55113
rect 12688 54915 12690 54971
rect 12690 54915 12742 54971
rect 12742 54915 12744 54971
rect 12688 54773 12690 54829
rect 12690 54773 12742 54829
rect 12742 54773 12744 54829
rect 12688 54631 12690 54687
rect 12690 54631 12742 54687
rect 12742 54631 12744 54687
rect 11350 54475 11352 54519
rect 11352 54475 11404 54519
rect 11404 54475 11406 54519
rect 11350 54463 11406 54475
rect 1896 53031 1952 53087
rect 1896 52889 1952 52945
rect 1896 52747 1952 52803
rect 1896 52605 1952 52661
rect 6106 53758 6108 53814
rect 6108 53758 6160 53814
rect 6160 53758 6162 53814
rect 4768 53673 4824 53729
rect 4768 53531 4770 53587
rect 4770 53531 4822 53587
rect 4822 53531 4824 53587
rect 4768 53389 4770 53445
rect 4770 53389 4822 53445
rect 4822 53389 4824 53445
rect 4768 53247 4770 53303
rect 4770 53247 4822 53303
rect 4822 53247 4824 53303
rect 4768 53105 4770 53161
rect 4770 53105 4822 53161
rect 4822 53105 4824 53161
rect 4768 52963 4824 53019
rect 4948 53673 5004 53729
rect 4948 53531 4950 53587
rect 4950 53531 5002 53587
rect 5002 53531 5004 53587
rect 4948 53389 4950 53445
rect 4950 53389 5002 53445
rect 5002 53389 5004 53445
rect 4948 53247 4950 53303
rect 4950 53247 5002 53303
rect 5002 53247 5004 53303
rect 4948 53105 4950 53161
rect 4950 53105 5002 53161
rect 5002 53105 5004 53161
rect 4948 52963 5004 53019
rect 5436 53673 5492 53729
rect 5436 53531 5438 53587
rect 5438 53531 5490 53587
rect 5490 53531 5492 53587
rect 5436 53389 5438 53445
rect 5438 53389 5490 53445
rect 5490 53389 5492 53445
rect 5436 53247 5438 53303
rect 5438 53247 5490 53303
rect 5490 53247 5492 53303
rect 5436 53105 5438 53161
rect 5438 53105 5490 53161
rect 5490 53105 5492 53161
rect 5436 52963 5492 53019
rect 5924 53673 5980 53729
rect 5924 53531 5926 53587
rect 5926 53531 5978 53587
rect 5978 53531 5980 53587
rect 5924 53389 5926 53445
rect 5926 53389 5978 53445
rect 5978 53389 5980 53445
rect 5924 53247 5926 53303
rect 5926 53247 5978 53303
rect 5978 53247 5980 53303
rect 5924 53105 5926 53161
rect 5926 53105 5978 53161
rect 5978 53105 5980 53161
rect 5924 52963 5980 53019
rect 6106 53616 6108 53672
rect 6108 53616 6160 53672
rect 6160 53616 6162 53672
rect 6106 53474 6108 53530
rect 6108 53474 6160 53530
rect 6160 53474 6162 53530
rect 6106 53332 6108 53388
rect 6108 53332 6160 53388
rect 6160 53332 6162 53388
rect 6106 53190 6108 53246
rect 6108 53190 6160 53246
rect 6160 53190 6162 53246
rect 6106 53048 6108 53104
rect 6108 53048 6160 53104
rect 6160 53048 6162 53104
rect 6106 52906 6162 52962
rect 6288 53673 6344 53729
rect 6288 53531 6290 53587
rect 6290 53531 6342 53587
rect 6342 53531 6344 53587
rect 6288 53389 6290 53445
rect 6290 53389 6342 53445
rect 6342 53389 6344 53445
rect 6288 53247 6290 53303
rect 6290 53247 6342 53303
rect 6342 53247 6344 53303
rect 6288 53105 6290 53161
rect 6290 53105 6342 53161
rect 6342 53105 6344 53161
rect 6288 52963 6344 53019
rect 6776 53673 6832 53729
rect 6776 53531 6778 53587
rect 6778 53531 6830 53587
rect 6830 53531 6832 53587
rect 6776 53389 6778 53445
rect 6778 53389 6830 53445
rect 6830 53389 6832 53445
rect 6776 53247 6778 53303
rect 6778 53247 6830 53303
rect 6830 53247 6832 53303
rect 6776 53105 6778 53161
rect 6778 53105 6830 53161
rect 6830 53105 6832 53161
rect 6776 52963 6832 53019
rect 1896 52463 1952 52519
rect 7264 53673 7320 53729
rect 7264 53531 7266 53587
rect 7266 53531 7318 53587
rect 7318 53531 7320 53587
rect 7264 53389 7266 53445
rect 7266 53389 7318 53445
rect 7318 53389 7320 53445
rect 7264 53247 7266 53303
rect 7266 53247 7318 53303
rect 7318 53247 7320 53303
rect 7264 53105 7266 53161
rect 7266 53105 7318 53161
rect 7318 53105 7320 53161
rect 7264 52963 7320 53019
rect 7444 53673 7500 53729
rect 7444 53531 7446 53587
rect 7446 53531 7498 53587
rect 7498 53531 7500 53587
rect 7444 53389 7446 53445
rect 7446 53389 7498 53445
rect 7498 53389 7500 53445
rect 7444 53247 7446 53303
rect 7446 53247 7498 53303
rect 7498 53247 7500 53303
rect 7444 53105 7446 53161
rect 7446 53105 7498 53161
rect 7498 53105 7500 53161
rect 7444 52963 7500 53019
rect 9179 53741 9235 53797
rect 9321 53741 9377 53797
rect 9463 53741 9519 53797
rect 11350 53758 11352 53814
rect 11352 53758 11404 53814
rect 11404 53758 11406 53814
rect 9179 53599 9235 53655
rect 9321 53599 9377 53655
rect 9463 53599 9519 53655
rect 9179 53457 9235 53513
rect 9321 53457 9377 53513
rect 9463 53457 9519 53513
rect 9179 53315 9235 53371
rect 9321 53315 9377 53371
rect 9463 53315 9519 53371
rect 9179 53173 9235 53229
rect 9321 53173 9377 53229
rect 9463 53173 9519 53229
rect 9179 53031 9235 53087
rect 9321 53031 9377 53087
rect 9463 53031 9519 53087
rect 10012 53673 10068 53729
rect 10012 53531 10014 53587
rect 10014 53531 10066 53587
rect 10066 53531 10068 53587
rect 10012 53389 10014 53445
rect 10014 53389 10066 53445
rect 10066 53389 10068 53445
rect 10012 53247 10014 53303
rect 10014 53247 10066 53303
rect 10066 53247 10068 53303
rect 10012 53105 10014 53161
rect 10014 53105 10066 53161
rect 10066 53105 10068 53161
rect 10012 52963 10068 53019
rect 10192 53673 10248 53729
rect 10192 53531 10194 53587
rect 10194 53531 10246 53587
rect 10246 53531 10248 53587
rect 10192 53389 10194 53445
rect 10194 53389 10246 53445
rect 10246 53389 10248 53445
rect 10192 53247 10194 53303
rect 10194 53247 10246 53303
rect 10246 53247 10248 53303
rect 10192 53105 10194 53161
rect 10194 53105 10246 53161
rect 10246 53105 10248 53161
rect 10192 52963 10248 53019
rect 10680 53673 10736 53729
rect 10680 53531 10682 53587
rect 10682 53531 10734 53587
rect 10734 53531 10736 53587
rect 10680 53389 10682 53445
rect 10682 53389 10734 53445
rect 10734 53389 10736 53445
rect 10680 53247 10682 53303
rect 10682 53247 10734 53303
rect 10734 53247 10736 53303
rect 10680 53105 10682 53161
rect 10682 53105 10734 53161
rect 10734 53105 10736 53161
rect 10680 52963 10736 53019
rect 11168 53673 11224 53729
rect 11168 53531 11170 53587
rect 11170 53531 11222 53587
rect 11222 53531 11224 53587
rect 11168 53389 11170 53445
rect 11170 53389 11222 53445
rect 11222 53389 11224 53445
rect 11168 53247 11170 53303
rect 11170 53247 11222 53303
rect 11222 53247 11224 53303
rect 11168 53105 11170 53161
rect 11170 53105 11222 53161
rect 11222 53105 11224 53161
rect 11168 52963 11224 53019
rect 11350 53616 11352 53672
rect 11352 53616 11404 53672
rect 11404 53616 11406 53672
rect 11350 53474 11352 53530
rect 11352 53474 11404 53530
rect 11404 53474 11406 53530
rect 11350 53332 11352 53388
rect 11352 53332 11404 53388
rect 11404 53332 11406 53388
rect 11350 53190 11352 53246
rect 11352 53190 11404 53246
rect 11404 53190 11406 53246
rect 11350 53048 11352 53104
rect 11352 53048 11404 53104
rect 11404 53048 11406 53104
rect 9179 52889 9235 52945
rect 9321 52889 9377 52945
rect 9463 52889 9519 52945
rect 11350 52906 11406 52962
rect 11532 53673 11588 53729
rect 11532 53531 11534 53587
rect 11534 53531 11586 53587
rect 11586 53531 11588 53587
rect 11532 53389 11534 53445
rect 11534 53389 11586 53445
rect 11586 53389 11588 53445
rect 11532 53247 11534 53303
rect 11534 53247 11586 53303
rect 11586 53247 11588 53303
rect 11532 53105 11534 53161
rect 11534 53105 11586 53161
rect 11586 53105 11588 53161
rect 11532 52963 11588 53019
rect 12020 53673 12076 53729
rect 12020 53531 12022 53587
rect 12022 53531 12074 53587
rect 12074 53531 12076 53587
rect 12020 53389 12022 53445
rect 12022 53389 12074 53445
rect 12074 53389 12076 53445
rect 12020 53247 12022 53303
rect 12022 53247 12074 53303
rect 12074 53247 12076 53303
rect 12020 53105 12022 53161
rect 12022 53105 12074 53161
rect 12074 53105 12076 53161
rect 12020 52963 12076 53019
rect 12508 53673 12564 53729
rect 12508 53531 12510 53587
rect 12510 53531 12562 53587
rect 12562 53531 12564 53587
rect 12508 53389 12510 53445
rect 12510 53389 12562 53445
rect 12562 53389 12564 53445
rect 12508 53247 12510 53303
rect 12510 53247 12562 53303
rect 12562 53247 12564 53303
rect 12508 53105 12510 53161
rect 12510 53105 12562 53161
rect 12562 53105 12564 53161
rect 12508 52963 12564 53019
rect 12688 53673 12744 53729
rect 12688 53531 12690 53587
rect 12690 53531 12742 53587
rect 12742 53531 12744 53587
rect 12688 53389 12690 53445
rect 12690 53389 12742 53445
rect 12742 53389 12744 53445
rect 12688 53247 12690 53303
rect 12690 53247 12742 53303
rect 12742 53247 12744 53303
rect 12688 53105 12690 53161
rect 12690 53105 12742 53161
rect 12742 53105 12744 53161
rect 12688 52963 12744 53019
rect 9179 52747 9235 52803
rect 9321 52747 9377 52803
rect 9463 52747 9519 52803
rect 9179 52605 9235 52661
rect 9321 52605 9377 52661
rect 9463 52605 9519 52661
rect 9179 52463 9235 52519
rect 9321 52463 9377 52519
rect 9463 52463 9519 52519
rect 3988 48916 4044 48918
rect 3988 48864 3990 48916
rect 3990 48864 4042 48916
rect 4042 48864 4044 48916
rect 3988 48862 4044 48864
rect 4112 48916 4168 48918
rect 4112 48864 4114 48916
rect 4114 48864 4166 48916
rect 4166 48864 4168 48916
rect 4112 48862 4168 48864
rect 4236 48916 4292 48918
rect 4236 48864 4238 48916
rect 4238 48864 4290 48916
rect 4290 48864 4292 48916
rect 4236 48862 4292 48864
rect 3988 48792 4044 48794
rect 3988 48740 3990 48792
rect 3990 48740 4042 48792
rect 4042 48740 4044 48792
rect 3988 48738 4044 48740
rect 4112 48792 4168 48794
rect 4112 48740 4114 48792
rect 4114 48740 4166 48792
rect 4166 48740 4168 48792
rect 4112 48738 4168 48740
rect 4236 48792 4292 48794
rect 4236 48740 4238 48792
rect 4238 48740 4290 48792
rect 4290 48740 4292 48792
rect 4236 48738 4292 48740
rect 3988 48668 4044 48670
rect 3988 48616 3990 48668
rect 3990 48616 4042 48668
rect 4042 48616 4044 48668
rect 3988 48614 4044 48616
rect 4112 48668 4168 48670
rect 4112 48616 4114 48668
rect 4114 48616 4166 48668
rect 4166 48616 4168 48668
rect 4112 48614 4168 48616
rect 4236 48668 4292 48670
rect 4236 48616 4238 48668
rect 4238 48616 4290 48668
rect 4290 48616 4292 48668
rect 4236 48614 4292 48616
rect 3988 48544 4044 48546
rect 3988 48492 3990 48544
rect 3990 48492 4042 48544
rect 4042 48492 4044 48544
rect 3988 48490 4044 48492
rect 4112 48544 4168 48546
rect 4112 48492 4114 48544
rect 4114 48492 4166 48544
rect 4166 48492 4168 48544
rect 4112 48490 4168 48492
rect 4236 48544 4292 48546
rect 4236 48492 4238 48544
rect 4238 48492 4290 48544
rect 4290 48492 4292 48544
rect 4236 48490 4292 48492
rect 3988 48420 4044 48422
rect 3988 48368 3990 48420
rect 3990 48368 4042 48420
rect 4042 48368 4044 48420
rect 3988 48366 4044 48368
rect 4112 48420 4168 48422
rect 4112 48368 4114 48420
rect 4114 48368 4166 48420
rect 4166 48368 4168 48420
rect 4112 48366 4168 48368
rect 4236 48420 4292 48422
rect 4236 48368 4238 48420
rect 4238 48368 4290 48420
rect 4290 48368 4292 48420
rect 4236 48366 4292 48368
rect 3988 48296 4044 48298
rect 3988 48244 3990 48296
rect 3990 48244 4042 48296
rect 4042 48244 4044 48296
rect 3988 48242 4044 48244
rect 4112 48296 4168 48298
rect 4112 48244 4114 48296
rect 4114 48244 4166 48296
rect 4166 48244 4168 48296
rect 4112 48242 4168 48244
rect 4236 48296 4292 48298
rect 4236 48244 4238 48296
rect 4238 48244 4290 48296
rect 4290 48244 4292 48296
rect 4236 48242 4292 48244
rect 3988 48172 4044 48174
rect 3988 48120 3990 48172
rect 3990 48120 4042 48172
rect 4042 48120 4044 48172
rect 3988 48118 4044 48120
rect 4112 48172 4168 48174
rect 4112 48120 4114 48172
rect 4114 48120 4166 48172
rect 4166 48120 4168 48172
rect 4112 48118 4168 48120
rect 4236 48172 4292 48174
rect 4236 48120 4238 48172
rect 4238 48120 4290 48172
rect 4290 48120 4292 48172
rect 4236 48118 4292 48120
rect 3988 48048 4044 48050
rect 3988 47996 3990 48048
rect 3990 47996 4042 48048
rect 4042 47996 4044 48048
rect 3988 47994 4044 47996
rect 4112 48048 4168 48050
rect 4112 47996 4114 48048
rect 4114 47996 4166 48048
rect 4166 47996 4168 48048
rect 4112 47994 4168 47996
rect 4236 48048 4292 48050
rect 4236 47996 4238 48048
rect 4238 47996 4290 48048
rect 4290 47996 4292 48048
rect 4236 47994 4292 47996
rect 3988 47924 4044 47926
rect 3988 47872 3990 47924
rect 3990 47872 4042 47924
rect 4042 47872 4044 47924
rect 3988 47870 4044 47872
rect 4112 47924 4168 47926
rect 4112 47872 4114 47924
rect 4114 47872 4166 47924
rect 4166 47872 4168 47924
rect 4112 47870 4168 47872
rect 4236 47924 4292 47926
rect 4236 47872 4238 47924
rect 4238 47872 4290 47924
rect 4290 47872 4292 47924
rect 4236 47870 4292 47872
rect 3988 47800 4044 47802
rect 3988 47748 3990 47800
rect 3990 47748 4042 47800
rect 4042 47748 4044 47800
rect 3988 47746 4044 47748
rect 4112 47800 4168 47802
rect 4112 47748 4114 47800
rect 4114 47748 4166 47800
rect 4166 47748 4168 47800
rect 4112 47746 4168 47748
rect 4236 47800 4292 47802
rect 4236 47748 4238 47800
rect 4238 47748 4290 47800
rect 4290 47748 4292 47800
rect 4236 47746 4292 47748
rect 3618 47358 3620 47414
rect 3620 47358 3672 47414
rect 3672 47358 3674 47414
rect 3618 47216 3620 47272
rect 3620 47216 3672 47272
rect 3672 47216 3674 47272
rect 3618 47074 3620 47130
rect 3620 47074 3672 47130
rect 3672 47074 3674 47130
rect 3618 46932 3620 46988
rect 3620 46932 3672 46988
rect 3672 46932 3674 46988
rect 3618 46790 3620 46846
rect 3620 46790 3672 46846
rect 3672 46790 3674 46846
rect 3618 46648 3620 46704
rect 3620 46648 3672 46704
rect 3672 46648 3674 46704
rect 3618 46506 3620 46562
rect 3620 46506 3672 46562
rect 3672 46506 3674 46562
rect 3618 46364 3620 46420
rect 3620 46364 3672 46420
rect 3672 46364 3674 46420
rect 11562 49512 11618 49568
rect 11674 49512 11730 49568
rect 11562 49400 11618 49456
rect 11674 49400 11730 49456
rect 11562 49288 11618 49344
rect 11674 49288 11730 49344
rect 10792 48990 10848 49014
rect 10792 48958 10794 48990
rect 10794 48958 10846 48990
rect 10846 48958 10848 48990
rect 10792 48816 10794 48872
rect 10794 48816 10846 48872
rect 10846 48816 10848 48872
rect 10792 48674 10794 48730
rect 10794 48674 10846 48730
rect 10846 48674 10848 48730
rect 10792 48532 10794 48588
rect 10794 48532 10846 48588
rect 10846 48532 10848 48588
rect 10792 48390 10794 48446
rect 10794 48390 10846 48446
rect 10846 48390 10848 48446
rect 10792 48248 10794 48304
rect 10794 48248 10846 48304
rect 10846 48248 10848 48304
rect 10792 48106 10794 48162
rect 10794 48106 10846 48162
rect 10846 48106 10848 48162
rect 10792 48002 10794 48020
rect 10794 48002 10846 48020
rect 10846 48002 10848 48020
rect 10792 47964 10848 48002
rect 11011 47341 11013 47397
rect 11013 47341 11065 47397
rect 11065 47341 11067 47397
rect 11011 47199 11013 47255
rect 11013 47199 11065 47255
rect 11065 47199 11067 47255
rect 11011 47057 11013 47113
rect 11013 47057 11065 47113
rect 11065 47057 11067 47113
rect 11011 46915 11013 46971
rect 11013 46915 11065 46971
rect 11065 46915 11067 46971
rect 11011 46773 11013 46829
rect 11013 46773 11065 46829
rect 11065 46773 11067 46829
rect 11011 46631 11013 46687
rect 11013 46631 11065 46687
rect 11065 46631 11067 46687
rect 3979 45339 4035 45341
rect 3979 45287 3981 45339
rect 3981 45287 4033 45339
rect 4033 45287 4035 45339
rect 3979 45285 4035 45287
rect 4103 45339 4159 45341
rect 4103 45287 4105 45339
rect 4105 45287 4157 45339
rect 4157 45287 4159 45339
rect 4103 45285 4159 45287
rect 4227 45339 4283 45341
rect 4227 45287 4229 45339
rect 4229 45287 4281 45339
rect 4281 45287 4283 45339
rect 4227 45285 4283 45287
rect 3979 45215 4035 45217
rect 3979 45163 3981 45215
rect 3981 45163 4033 45215
rect 4033 45163 4035 45215
rect 3979 45161 4035 45163
rect 4103 45215 4159 45217
rect 4103 45163 4105 45215
rect 4105 45163 4157 45215
rect 4157 45163 4159 45215
rect 4103 45161 4159 45163
rect 4227 45215 4283 45217
rect 4227 45163 4229 45215
rect 4229 45163 4281 45215
rect 4281 45163 4283 45215
rect 4227 45161 4283 45163
rect 3979 45091 4035 45093
rect 3979 45039 3981 45091
rect 3981 45039 4033 45091
rect 4033 45039 4035 45091
rect 3979 45037 4035 45039
rect 4103 45091 4159 45093
rect 4103 45039 4105 45091
rect 4105 45039 4157 45091
rect 4157 45039 4159 45091
rect 4103 45037 4159 45039
rect 4227 45091 4283 45093
rect 4227 45039 4229 45091
rect 4229 45039 4281 45091
rect 4281 45039 4283 45091
rect 4227 45037 4283 45039
rect 3979 44967 4035 44969
rect 3979 44915 3981 44967
rect 3981 44915 4033 44967
rect 4033 44915 4035 44967
rect 3979 44913 4035 44915
rect 4103 44967 4159 44969
rect 4103 44915 4105 44967
rect 4105 44915 4157 44967
rect 4157 44915 4159 44967
rect 4103 44913 4159 44915
rect 4227 44967 4283 44969
rect 4227 44915 4229 44967
rect 4229 44915 4281 44967
rect 4281 44915 4283 44967
rect 4227 44913 4283 44915
rect 3979 44843 4035 44845
rect 3979 44791 3981 44843
rect 3981 44791 4033 44843
rect 4033 44791 4035 44843
rect 3979 44789 4035 44791
rect 4103 44843 4159 44845
rect 4103 44791 4105 44843
rect 4105 44791 4157 44843
rect 4157 44791 4159 44843
rect 4103 44789 4159 44791
rect 4227 44843 4283 44845
rect 4227 44791 4229 44843
rect 4229 44791 4281 44843
rect 4281 44791 4283 44843
rect 4227 44789 4283 44791
rect 3979 44719 4035 44721
rect 3979 44667 3981 44719
rect 3981 44667 4033 44719
rect 4033 44667 4035 44719
rect 3979 44665 4035 44667
rect 4103 44719 4159 44721
rect 4103 44667 4105 44719
rect 4105 44667 4157 44719
rect 4157 44667 4159 44719
rect 4103 44665 4159 44667
rect 4227 44719 4283 44721
rect 4227 44667 4229 44719
rect 4229 44667 4281 44719
rect 4281 44667 4283 44719
rect 4227 44665 4283 44667
rect 3979 44595 4035 44597
rect 3979 44543 3981 44595
rect 3981 44543 4033 44595
rect 4033 44543 4035 44595
rect 3979 44541 4035 44543
rect 4103 44595 4159 44597
rect 4103 44543 4105 44595
rect 4105 44543 4157 44595
rect 4157 44543 4159 44595
rect 4103 44541 4159 44543
rect 4227 44595 4283 44597
rect 4227 44543 4229 44595
rect 4229 44543 4281 44595
rect 4281 44543 4283 44595
rect 4227 44541 4283 44543
rect 3618 44180 3674 44197
rect 3618 44141 3620 44180
rect 3620 44141 3672 44180
rect 3672 44141 3674 44180
rect 3618 43999 3620 44055
rect 3620 43999 3672 44055
rect 3672 43999 3674 44055
rect 3618 43857 3620 43913
rect 3620 43857 3672 43913
rect 3672 43857 3674 43913
rect 3618 43715 3620 43771
rect 3620 43715 3672 43771
rect 3672 43715 3674 43771
rect 3618 43573 3620 43629
rect 3620 43573 3672 43629
rect 3672 43573 3674 43629
rect 3618 43431 3620 43487
rect 3620 43431 3672 43487
rect 3672 43431 3674 43487
rect 3618 43289 3620 43345
rect 3620 43289 3672 43345
rect 3672 43289 3674 43345
rect 3618 43147 3620 43203
rect 3620 43147 3672 43203
rect 3672 43147 3674 43203
rect 3618 43005 3620 43061
rect 3620 43005 3672 43061
rect 3672 43005 3674 43061
rect 3618 42880 3620 42919
rect 3620 42880 3672 42919
rect 3672 42880 3674 42919
rect 3618 42863 3674 42880
rect 3618 42580 3674 42597
rect 3618 42541 3620 42580
rect 3620 42541 3672 42580
rect 3672 42541 3674 42580
rect 3618 42399 3620 42455
rect 3620 42399 3672 42455
rect 3672 42399 3674 42455
rect 3618 42257 3620 42313
rect 3620 42257 3672 42313
rect 3672 42257 3674 42313
rect 3618 42115 3620 42171
rect 3620 42115 3672 42171
rect 3672 42115 3674 42171
rect 3618 41973 3620 42029
rect 3620 41973 3672 42029
rect 3672 41973 3674 42029
rect 3618 41831 3620 41887
rect 3620 41831 3672 41887
rect 3672 41831 3674 41887
rect 3618 41689 3620 41745
rect 3620 41689 3672 41745
rect 3672 41689 3674 41745
rect 3618 41547 3620 41603
rect 3620 41547 3672 41603
rect 3672 41547 3674 41603
rect 3618 41405 3620 41461
rect 3620 41405 3672 41461
rect 3672 41405 3674 41461
rect 3618 41280 3620 41319
rect 3620 41280 3672 41319
rect 3672 41280 3674 41319
rect 3618 41263 3674 41280
rect 1846 40700 1902 40702
rect 1988 40700 2044 40702
rect 2130 40700 2186 40702
rect 2272 40700 2328 40702
rect 2414 40700 2470 40702
rect 2556 40700 2612 40702
rect 2698 40700 2754 40702
rect 2840 40700 2896 40702
rect 2982 40700 3038 40702
rect 3124 40700 3180 40702
rect 3266 40700 3322 40702
rect 3408 40700 3464 40702
rect 3550 40700 3606 40702
rect 1846 40648 1848 40700
rect 1848 40648 1902 40700
rect 1988 40648 2044 40700
rect 2130 40648 2186 40700
rect 2272 40648 2328 40700
rect 2414 40648 2470 40700
rect 2556 40648 2612 40700
rect 2698 40648 2754 40700
rect 2840 40648 2896 40700
rect 2982 40648 3038 40700
rect 3124 40648 3180 40700
rect 3266 40648 3322 40700
rect 3408 40648 3464 40700
rect 3550 40648 3606 40700
rect 1846 40646 1902 40648
rect 1988 40646 2044 40648
rect 2130 40646 2186 40648
rect 2272 40646 2328 40648
rect 2414 40646 2470 40648
rect 2556 40646 2612 40648
rect 2698 40646 2754 40648
rect 2840 40646 2896 40648
rect 2982 40646 3038 40648
rect 3124 40646 3180 40648
rect 3266 40646 3322 40648
rect 3408 40646 3464 40648
rect 3550 40646 3606 40648
rect 3692 40646 3748 40702
rect 1781 39418 1837 39420
rect 1781 39364 1783 39418
rect 1783 39364 1835 39418
rect 1835 39364 1837 39418
rect 1781 39222 1783 39278
rect 1783 39222 1835 39278
rect 1835 39222 1837 39278
rect 1781 39080 1783 39136
rect 1783 39080 1835 39136
rect 1835 39080 1837 39136
rect 1781 38938 1783 38994
rect 1783 38938 1835 38994
rect 1835 38938 1837 38994
rect 1781 38846 1783 38852
rect 1783 38846 1835 38852
rect 1835 38846 1837 38852
rect 1781 38796 1837 38846
rect 2438 39944 2494 39946
rect 2580 39944 2636 39946
rect 2722 39944 2778 39946
rect 2864 39944 2920 39946
rect 3006 39944 3062 39946
rect 3148 39944 3204 39946
rect 3290 39944 3346 39946
rect 3432 39944 3488 39946
rect 3574 39944 3630 39946
rect 3716 39944 3772 39946
rect 3858 39944 3914 39946
rect 4000 39944 4056 39946
rect 4142 39944 4198 39946
rect 4284 39944 4340 39946
rect 4426 39944 4482 39946
rect 2438 39892 2445 39944
rect 2445 39892 2494 39944
rect 2580 39892 2636 39944
rect 2722 39892 2778 39944
rect 2864 39892 2920 39944
rect 3006 39892 3062 39944
rect 3148 39892 3204 39944
rect 3290 39892 3346 39944
rect 3432 39892 3488 39944
rect 3574 39892 3630 39944
rect 3716 39892 3772 39944
rect 3858 39892 3914 39944
rect 4000 39892 4056 39944
rect 4142 39892 4198 39944
rect 4284 39892 4340 39944
rect 4426 39892 4473 39944
rect 4473 39892 4482 39944
rect 2438 39890 2494 39892
rect 2580 39890 2636 39892
rect 2722 39890 2778 39892
rect 2864 39890 2920 39892
rect 3006 39890 3062 39892
rect 3148 39890 3204 39892
rect 3290 39890 3346 39892
rect 3432 39890 3488 39892
rect 3574 39890 3630 39892
rect 3716 39890 3772 39892
rect 3858 39890 3914 39892
rect 4000 39890 4056 39892
rect 4142 39890 4198 39892
rect 4284 39890 4340 39892
rect 4426 39890 4482 39892
rect 5093 39418 5149 39420
rect 5093 39364 5095 39418
rect 5095 39364 5147 39418
rect 5147 39364 5149 39418
rect 5093 39222 5095 39278
rect 5095 39222 5147 39278
rect 5147 39222 5149 39278
rect 5093 39080 5095 39136
rect 5095 39080 5147 39136
rect 5147 39080 5149 39136
rect 5093 38938 5095 38994
rect 5095 38938 5147 38994
rect 5147 38938 5149 38994
rect 5093 38846 5095 38852
rect 5095 38846 5147 38852
rect 5147 38846 5149 38852
rect 5093 38796 5149 38846
rect 6059 39358 6061 39414
rect 6061 39358 6113 39414
rect 6113 39358 6115 39414
rect 6059 39216 6061 39272
rect 6061 39216 6113 39272
rect 6113 39216 6115 39272
rect 6059 39074 6061 39130
rect 6061 39074 6113 39130
rect 6113 39074 6115 39130
rect 6059 38932 6061 38988
rect 6061 38932 6113 38988
rect 6113 38932 6115 38988
rect 6059 38790 6061 38846
rect 6061 38790 6113 38846
rect 6113 38790 6115 38846
rect 7025 39418 7081 39420
rect 7025 39364 7027 39418
rect 7027 39364 7079 39418
rect 7079 39364 7081 39418
rect 7025 39222 7027 39278
rect 7027 39222 7079 39278
rect 7079 39222 7081 39278
rect 7025 39080 7027 39136
rect 7027 39080 7079 39136
rect 7079 39080 7081 39136
rect 7025 38938 7027 38994
rect 7027 38938 7079 38994
rect 7079 38938 7081 38994
rect 7025 38846 7027 38852
rect 7027 38846 7079 38852
rect 7079 38846 7081 38852
rect 7025 38796 7081 38846
rect 6059 38648 6061 38704
rect 6061 38648 6113 38704
rect 6113 38648 6115 38704
rect 6059 38506 6061 38562
rect 6061 38506 6113 38562
rect 6113 38506 6115 38562
rect 6059 38364 6115 38420
rect 56 37780 112 37797
rect 56 37741 58 37780
rect 58 37741 110 37780
rect 110 37741 112 37780
rect 56 37599 58 37655
rect 58 37599 110 37655
rect 110 37599 112 37655
rect 56 37457 58 37513
rect 58 37457 110 37513
rect 110 37457 112 37513
rect 56 37315 58 37371
rect 58 37315 110 37371
rect 110 37315 112 37371
rect 56 37173 58 37229
rect 58 37173 110 37229
rect 110 37173 112 37229
rect 56 37031 58 37087
rect 58 37031 110 37087
rect 110 37031 112 37087
rect 56 36889 58 36945
rect 58 36889 110 36945
rect 110 36889 112 36945
rect 56 36747 58 36803
rect 58 36747 110 36803
rect 110 36747 112 36803
rect 56 36605 58 36661
rect 58 36605 110 36661
rect 110 36605 112 36661
rect 56 36480 58 36519
rect 58 36480 110 36519
rect 110 36480 112 36519
rect 56 36463 112 36480
rect 734 37741 790 37797
rect 734 37599 790 37655
rect 734 37457 790 37513
rect 734 37315 790 37371
rect 734 37173 790 37229
rect 876 37741 932 37797
rect 1018 37741 1074 37797
rect 876 37599 932 37655
rect 1018 37599 1074 37655
rect 876 37457 932 37513
rect 1018 37457 1074 37513
rect 876 37315 932 37371
rect 1018 37315 1074 37371
rect 876 37173 932 37229
rect 1018 37173 1074 37229
rect 734 37031 790 37087
rect 876 37031 932 37087
rect 1018 37031 1074 37087
rect 734 36889 790 36945
rect 876 36889 932 36945
rect 1018 36889 1074 36945
rect 734 36747 790 36803
rect 876 36747 932 36803
rect 1018 36747 1074 36803
rect 734 36605 790 36661
rect 876 36605 932 36661
rect 1018 36605 1074 36661
rect 734 36463 790 36519
rect 876 36463 932 36519
rect 1018 36463 1074 36519
rect 175 36122 231 36178
rect 317 36122 373 36178
rect 175 35980 231 36036
rect 317 35980 373 36036
rect 175 35838 231 35894
rect 317 35838 373 35894
rect 175 35696 231 35752
rect 317 35696 373 35752
rect 175 35554 231 35610
rect 317 35554 373 35610
rect 175 35412 231 35468
rect 317 35412 373 35468
rect 175 35270 231 35326
rect 317 35270 373 35326
rect 175 35128 231 35184
rect 317 35128 373 35184
rect 175 34986 231 35042
rect 317 34986 373 35042
rect 175 34844 231 34900
rect 317 34844 373 34900
rect 175 34702 231 34758
rect 317 34702 373 34758
rect 175 34560 231 34616
rect 317 34560 373 34616
rect 175 34418 231 34474
rect 317 34418 373 34474
rect 175 34276 231 34332
rect 317 34276 373 34332
rect 175 34134 231 34190
rect 317 34134 373 34190
rect 175 33992 231 34048
rect 317 33992 373 34048
rect 175 33850 231 33906
rect 317 33850 373 33906
rect 175 33708 231 33764
rect 317 33708 373 33764
rect 496 35576 552 35617
rect 496 35561 498 35576
rect 498 35561 550 35576
rect 550 35561 552 35576
rect 496 35419 498 35475
rect 498 35419 550 35475
rect 550 35419 552 35475
rect 496 35277 498 35333
rect 498 35277 550 35333
rect 550 35277 552 35333
rect 496 35135 498 35191
rect 498 35135 550 35191
rect 550 35135 552 35191
rect 496 34993 498 35049
rect 498 34993 550 35049
rect 550 34993 552 35049
rect 496 34851 498 34907
rect 498 34851 550 34907
rect 550 34851 552 34907
rect 496 34709 498 34765
rect 498 34709 550 34765
rect 550 34709 552 34765
rect 496 34567 498 34623
rect 498 34567 550 34623
rect 550 34567 552 34623
rect 496 34425 498 34481
rect 498 34425 550 34481
rect 550 34425 552 34481
rect 496 34283 498 34339
rect 498 34283 550 34339
rect 550 34283 552 34339
rect 496 34141 498 34197
rect 498 34141 550 34197
rect 550 34141 552 34197
rect 734 35576 790 35612
rect 734 35556 736 35576
rect 736 35556 788 35576
rect 788 35556 790 35576
rect 734 35414 736 35470
rect 736 35414 788 35470
rect 788 35414 790 35470
rect 734 35272 736 35328
rect 736 35272 788 35328
rect 788 35272 790 35328
rect 734 35130 736 35186
rect 736 35130 788 35186
rect 788 35130 790 35186
rect 734 34988 736 35044
rect 736 34988 788 35044
rect 788 34988 790 35044
rect 734 34846 736 34902
rect 736 34846 788 34902
rect 788 34846 790 34902
rect 734 34704 736 34760
rect 736 34704 788 34760
rect 788 34704 790 34760
rect 734 34562 736 34618
rect 736 34562 788 34618
rect 788 34562 790 34618
rect 734 34420 736 34476
rect 736 34420 788 34476
rect 788 34420 790 34476
rect 734 34278 736 34334
rect 736 34278 788 34334
rect 788 34278 790 34334
rect 734 34172 736 34192
rect 736 34172 788 34192
rect 788 34172 790 34192
rect 734 34136 790 34172
rect 496 33999 498 34055
rect 498 33999 550 34055
rect 550 33999 552 34055
rect 496 33857 498 33913
rect 498 33857 550 33913
rect 550 33857 552 33913
rect 496 33756 498 33771
rect 498 33756 550 33771
rect 550 33756 552 33771
rect 496 33715 552 33756
rect 175 33566 231 33622
rect 317 33566 373 33622
rect 175 33424 231 33480
rect 317 33424 373 33480
rect 175 33282 231 33338
rect 317 33282 373 33338
rect 496 32922 498 32978
rect 498 32922 550 32978
rect 550 32922 552 32978
rect 496 32780 498 32836
rect 498 32780 550 32836
rect 550 32780 552 32836
rect 496 32638 498 32694
rect 498 32638 550 32694
rect 550 32638 552 32694
rect 496 32496 498 32552
rect 498 32496 550 32552
rect 550 32496 552 32552
rect 6059 37741 6061 37797
rect 6061 37741 6113 37797
rect 6113 37741 6115 37797
rect 6059 37599 6061 37655
rect 6061 37599 6113 37655
rect 6113 37599 6115 37655
rect 6059 37457 6061 37513
rect 6061 37457 6113 37513
rect 6113 37457 6115 37513
rect 6059 37315 6061 37371
rect 6061 37315 6113 37371
rect 6113 37315 6115 37371
rect 6059 37173 6061 37229
rect 6061 37173 6113 37229
rect 6113 37173 6115 37229
rect 6059 37031 6115 37087
rect 6059 36889 6115 36945
rect 6059 36747 6115 36803
rect 6059 36605 6115 36661
rect 6059 36463 6115 36519
rect 3102 35576 3158 35612
rect 3102 35556 3104 35576
rect 3104 35556 3156 35576
rect 3156 35556 3158 35576
rect 3102 35414 3104 35470
rect 3104 35414 3156 35470
rect 3156 35414 3158 35470
rect 3102 35272 3104 35328
rect 3104 35272 3156 35328
rect 3156 35272 3158 35328
rect 3102 35130 3104 35186
rect 3104 35130 3156 35186
rect 3156 35130 3158 35186
rect 3102 34988 3104 35044
rect 3104 34988 3156 35044
rect 3156 34988 3158 35044
rect 3102 34846 3104 34902
rect 3104 34846 3156 34902
rect 3156 34846 3158 34902
rect 3102 34704 3104 34760
rect 3104 34704 3156 34760
rect 3156 34704 3158 34760
rect 3102 34562 3104 34618
rect 3104 34562 3156 34618
rect 3156 34562 3158 34618
rect 3102 34420 3104 34476
rect 3104 34420 3156 34476
rect 3156 34420 3158 34476
rect 3102 34278 3104 34334
rect 3104 34278 3156 34334
rect 3156 34278 3158 34334
rect 3102 34172 3104 34192
rect 3104 34172 3156 34192
rect 3156 34172 3158 34192
rect 3102 34136 3158 34172
rect 4000 35660 4056 35716
rect 4000 35518 4002 35574
rect 4002 35518 4054 35574
rect 4054 35518 4056 35574
rect 4000 35376 4002 35432
rect 4002 35376 4054 35432
rect 4054 35376 4056 35432
rect 4000 35234 4002 35290
rect 4002 35234 4054 35290
rect 4054 35234 4056 35290
rect 4000 35092 4002 35148
rect 4002 35092 4054 35148
rect 4054 35092 4056 35148
rect 4000 34950 4002 35006
rect 4002 34950 4054 35006
rect 4054 34950 4056 35006
rect 4000 34808 4002 34864
rect 4002 34808 4054 34864
rect 4054 34808 4056 34864
rect 4000 34666 4002 34722
rect 4002 34666 4054 34722
rect 4054 34666 4056 34722
rect 4000 34524 4002 34580
rect 4002 34524 4054 34580
rect 4054 34524 4056 34580
rect 4000 34382 4002 34438
rect 4002 34382 4054 34438
rect 4054 34382 4056 34438
rect 4000 34240 4002 34296
rect 4002 34240 4054 34296
rect 4054 34240 4056 34296
rect 4000 34098 4002 34154
rect 4002 34098 4054 34154
rect 4054 34098 4056 34154
rect 4000 33956 4002 34012
rect 4002 33956 4054 34012
rect 4054 33956 4056 34012
rect 4898 35576 4954 35612
rect 4898 35556 4900 35576
rect 4900 35556 4952 35576
rect 4952 35556 4954 35576
rect 4898 35414 4900 35470
rect 4900 35414 4952 35470
rect 4952 35414 4954 35470
rect 4898 35272 4900 35328
rect 4900 35272 4952 35328
rect 4952 35272 4954 35328
rect 4898 35130 4900 35186
rect 4900 35130 4952 35186
rect 4952 35130 4954 35186
rect 4898 34988 4900 35044
rect 4900 34988 4952 35044
rect 4952 34988 4954 35044
rect 4898 34846 4900 34902
rect 4900 34846 4952 34902
rect 4952 34846 4954 34902
rect 4898 34704 4900 34760
rect 4900 34704 4952 34760
rect 4952 34704 4954 34760
rect 4898 34562 4900 34618
rect 4900 34562 4952 34618
rect 4952 34562 4954 34618
rect 4898 34420 4900 34476
rect 4900 34420 4952 34476
rect 4952 34420 4954 34476
rect 4898 34278 4900 34334
rect 4900 34278 4952 34334
rect 4952 34278 4954 34334
rect 4898 34172 4900 34192
rect 4900 34172 4952 34192
rect 4952 34172 4954 34192
rect 4898 34136 4954 34172
rect 4000 33814 4002 33870
rect 4002 33814 4054 33870
rect 4054 33814 4056 33870
rect 4000 33672 4002 33728
rect 4002 33672 4054 33728
rect 4054 33672 4056 33728
rect 4000 33530 4002 33586
rect 4002 33530 4054 33586
rect 4054 33530 4056 33586
rect 4000 33388 4002 33444
rect 4002 33388 4054 33444
rect 4054 33388 4056 33444
rect 4000 33246 4002 33302
rect 4002 33246 4054 33302
rect 4054 33246 4056 33302
rect 496 32354 498 32410
rect 498 32354 550 32410
rect 550 32354 552 32410
rect 4000 32479 4056 32535
rect 4000 32337 4002 32393
rect 4002 32337 4054 32393
rect 4054 32337 4056 32393
rect 496 32212 498 32268
rect 498 32212 550 32268
rect 550 32212 552 32268
rect 496 32070 498 32126
rect 498 32070 550 32126
rect 550 32070 552 32126
rect 496 31928 498 31984
rect 498 31928 550 31984
rect 550 31928 552 31984
rect 496 31786 498 31842
rect 498 31786 550 31842
rect 550 31786 552 31842
rect 496 31644 498 31700
rect 498 31644 550 31700
rect 550 31644 552 31700
rect 496 31502 498 31558
rect 498 31502 550 31558
rect 550 31502 552 31558
rect 496 31360 498 31416
rect 498 31360 550 31416
rect 550 31360 552 31416
rect 496 31218 498 31274
rect 498 31218 550 31274
rect 550 31218 552 31274
rect 496 31076 498 31132
rect 498 31076 550 31132
rect 550 31076 552 31132
rect 496 30934 498 30990
rect 498 30934 550 30990
rect 550 30934 552 30990
rect 496 30792 498 30848
rect 498 30792 550 30848
rect 550 30792 552 30848
rect 496 30650 498 30706
rect 498 30650 550 30706
rect 550 30650 552 30706
rect 496 30508 498 30564
rect 498 30508 550 30564
rect 550 30508 552 30564
rect 496 30366 498 30422
rect 498 30366 550 30422
rect 550 30366 552 30422
rect 496 30224 498 30280
rect 498 30224 550 30280
rect 550 30224 552 30280
rect 496 30082 498 30138
rect 498 30082 550 30138
rect 550 30082 552 30138
rect 978 32320 1034 32322
rect 978 32266 980 32320
rect 980 32266 1032 32320
rect 1032 32266 1034 32320
rect 978 32124 980 32180
rect 980 32124 1032 32180
rect 1032 32124 1034 32180
rect 978 31982 980 32038
rect 980 31982 1032 32038
rect 1032 31982 1034 32038
rect 978 31840 980 31896
rect 980 31840 1032 31896
rect 1032 31840 1034 31896
rect 978 31698 980 31754
rect 980 31698 1032 31754
rect 1032 31698 1034 31754
rect 978 31556 980 31612
rect 980 31556 1032 31612
rect 1032 31556 1034 31612
rect 978 31414 980 31470
rect 980 31414 1032 31470
rect 1032 31414 1034 31470
rect 978 31272 980 31328
rect 980 31272 1032 31328
rect 1032 31272 1034 31328
rect 978 31130 980 31186
rect 980 31130 1032 31186
rect 1032 31130 1034 31186
rect 978 30988 980 31044
rect 980 30988 1032 31044
rect 1032 30988 1034 31044
rect 978 30846 980 30902
rect 980 30846 1032 30902
rect 1032 30846 1034 30902
rect 978 30704 980 30760
rect 980 30704 1032 30760
rect 1032 30704 1034 30760
rect 978 30562 980 30618
rect 980 30562 1032 30618
rect 1032 30562 1034 30618
rect 978 30420 980 30476
rect 980 30420 1032 30476
rect 1032 30420 1034 30476
rect 978 30278 980 30334
rect 980 30278 1032 30334
rect 1032 30278 1034 30334
rect 2370 32320 2426 32322
rect 2370 32266 2372 32320
rect 2372 32266 2424 32320
rect 2424 32266 2426 32320
rect 2370 32124 2372 32180
rect 2372 32124 2424 32180
rect 2424 32124 2426 32180
rect 2370 31982 2372 32038
rect 2372 31982 2424 32038
rect 2424 31982 2426 32038
rect 2370 31840 2372 31896
rect 2372 31840 2424 31896
rect 2424 31840 2426 31896
rect 2370 31698 2372 31754
rect 2372 31698 2424 31754
rect 2424 31698 2426 31754
rect 2370 31556 2372 31612
rect 2372 31556 2424 31612
rect 2424 31556 2426 31612
rect 2370 31414 2372 31470
rect 2372 31414 2424 31470
rect 2424 31414 2426 31470
rect 2370 31272 2372 31328
rect 2372 31272 2424 31328
rect 2424 31272 2426 31328
rect 2370 31130 2372 31186
rect 2372 31130 2424 31186
rect 2424 31130 2426 31186
rect 2370 30988 2372 31044
rect 2372 30988 2424 31044
rect 2424 30988 2426 31044
rect 2370 30846 2372 30902
rect 2372 30846 2424 30902
rect 2424 30846 2426 30902
rect 2370 30704 2372 30760
rect 2372 30704 2424 30760
rect 2424 30704 2426 30760
rect 2370 30562 2372 30618
rect 2372 30562 2424 30618
rect 2424 30562 2426 30618
rect 2370 30420 2372 30476
rect 2372 30420 2424 30476
rect 2424 30420 2426 30476
rect 978 30136 980 30192
rect 980 30136 1032 30192
rect 1032 30136 1034 30192
rect 2370 30278 2372 30334
rect 2372 30278 2424 30334
rect 2424 30278 2426 30334
rect 2370 30136 2372 30192
rect 2372 30136 2424 30192
rect 2424 30136 2426 30192
rect 2786 32320 2842 32322
rect 2786 32266 2788 32320
rect 2788 32266 2840 32320
rect 2840 32266 2842 32320
rect 2786 32124 2788 32180
rect 2788 32124 2840 32180
rect 2840 32124 2842 32180
rect 2786 31982 2788 32038
rect 2788 31982 2840 32038
rect 2840 31982 2842 32038
rect 2786 31840 2788 31896
rect 2788 31840 2840 31896
rect 2840 31840 2842 31896
rect 2786 31698 2788 31754
rect 2788 31698 2840 31754
rect 2840 31698 2842 31754
rect 2786 31556 2788 31612
rect 2788 31556 2840 31612
rect 2840 31556 2842 31612
rect 2786 31414 2788 31470
rect 2788 31414 2840 31470
rect 2840 31414 2842 31470
rect 2786 31272 2788 31328
rect 2788 31272 2840 31328
rect 2840 31272 2842 31328
rect 2786 31130 2788 31186
rect 2788 31130 2840 31186
rect 2840 31130 2842 31186
rect 2786 30988 2788 31044
rect 2788 30988 2840 31044
rect 2840 30988 2842 31044
rect 2786 30846 2788 30902
rect 2788 30846 2840 30902
rect 2840 30846 2842 30902
rect 2786 30704 2788 30760
rect 2788 30704 2840 30760
rect 2840 30704 2842 30760
rect 3274 32320 3330 32323
rect 3274 32267 3276 32320
rect 3276 32267 3328 32320
rect 3328 32267 3330 32320
rect 3274 32125 3276 32181
rect 3276 32125 3328 32181
rect 3328 32125 3330 32181
rect 3274 31983 3276 32039
rect 3276 31983 3328 32039
rect 3328 31983 3330 32039
rect 3274 31841 3276 31897
rect 3276 31841 3328 31897
rect 3328 31841 3330 31897
rect 3274 31699 3276 31755
rect 3276 31699 3328 31755
rect 3328 31699 3330 31755
rect 3274 31557 3276 31613
rect 3276 31557 3328 31613
rect 3328 31557 3330 31613
rect 3274 31415 3276 31471
rect 3276 31415 3328 31471
rect 3328 31415 3330 31471
rect 3274 31273 3276 31329
rect 3276 31273 3328 31329
rect 3328 31273 3330 31329
rect 3274 31131 3276 31187
rect 3276 31131 3328 31187
rect 3328 31131 3330 31187
rect 3274 30989 3276 31045
rect 3276 30989 3328 31045
rect 3328 30989 3330 31045
rect 3274 30847 3276 30903
rect 3276 30847 3328 30903
rect 3328 30847 3330 30903
rect 3274 30708 3276 30761
rect 3276 30708 3328 30761
rect 3328 30708 3330 30761
rect 3274 30705 3330 30708
rect 3762 32270 3818 32272
rect 3762 32216 3764 32270
rect 3764 32216 3816 32270
rect 3816 32216 3818 32270
rect 3762 32074 3764 32130
rect 3764 32074 3816 32130
rect 3816 32074 3818 32130
rect 3762 31932 3764 31988
rect 3764 31932 3816 31988
rect 3816 31932 3818 31988
rect 3762 31790 3764 31846
rect 3764 31790 3816 31846
rect 3816 31790 3818 31846
rect 3762 31648 3764 31704
rect 3764 31648 3816 31704
rect 3816 31648 3818 31704
rect 3762 31506 3764 31562
rect 3764 31506 3816 31562
rect 3816 31506 3818 31562
rect 3762 31364 3764 31420
rect 3764 31364 3816 31420
rect 3816 31364 3818 31420
rect 3762 31222 3764 31278
rect 3764 31222 3816 31278
rect 3816 31222 3818 31278
rect 3762 31080 3764 31136
rect 3764 31080 3816 31136
rect 3816 31080 3818 31136
rect 3762 30938 3764 30994
rect 3764 30938 3816 30994
rect 3816 30938 3818 30994
rect 3762 30796 3764 30852
rect 3764 30796 3816 30852
rect 3816 30796 3818 30852
rect 3762 30658 3764 30710
rect 3764 30658 3816 30710
rect 3816 30658 3818 30710
rect 3762 30654 3818 30658
rect 4000 32195 4002 32251
rect 4002 32195 4054 32251
rect 4054 32195 4056 32251
rect 4000 32053 4002 32109
rect 4002 32053 4054 32109
rect 4054 32053 4056 32109
rect 4000 31911 4002 31967
rect 4002 31911 4054 31967
rect 4054 31911 4056 31967
rect 4000 31769 4002 31825
rect 4002 31769 4054 31825
rect 4054 31769 4056 31825
rect 4000 31627 4002 31683
rect 4002 31627 4054 31683
rect 4054 31627 4056 31683
rect 4000 31485 4002 31541
rect 4002 31485 4054 31541
rect 4054 31485 4056 31541
rect 4000 31343 4002 31399
rect 4002 31343 4054 31399
rect 4054 31343 4056 31399
rect 4000 31201 4002 31257
rect 4002 31201 4054 31257
rect 4054 31201 4056 31257
rect 4000 31059 4002 31115
rect 4002 31059 4054 31115
rect 4054 31059 4056 31115
rect 4000 30917 4002 30973
rect 4002 30917 4054 30973
rect 4054 30917 4056 30973
rect 4000 30775 4002 30831
rect 4002 30775 4054 30831
rect 4054 30775 4056 30831
rect 4000 30635 4002 30689
rect 4002 30635 4054 30689
rect 4054 30635 4056 30689
rect 4000 30633 4056 30635
rect 4238 32270 4294 32272
rect 4238 32216 4240 32270
rect 4240 32216 4292 32270
rect 4292 32216 4294 32270
rect 4238 32074 4240 32130
rect 4240 32074 4292 32130
rect 4292 32074 4294 32130
rect 4238 31932 4240 31988
rect 4240 31932 4292 31988
rect 4292 31932 4294 31988
rect 4238 31790 4240 31846
rect 4240 31790 4292 31846
rect 4292 31790 4294 31846
rect 4238 31648 4240 31704
rect 4240 31648 4292 31704
rect 4292 31648 4294 31704
rect 4238 31506 4240 31562
rect 4240 31506 4292 31562
rect 4292 31506 4294 31562
rect 4238 31364 4240 31420
rect 4240 31364 4292 31420
rect 4292 31364 4294 31420
rect 4238 31222 4240 31278
rect 4240 31222 4292 31278
rect 4292 31222 4294 31278
rect 4238 31080 4240 31136
rect 4240 31080 4292 31136
rect 4292 31080 4294 31136
rect 4238 30938 4240 30994
rect 4240 30938 4292 30994
rect 4292 30938 4294 30994
rect 4238 30796 4240 30852
rect 4240 30796 4292 30852
rect 4292 30796 4294 30852
rect 4238 30658 4240 30710
rect 4240 30658 4292 30710
rect 4292 30658 4294 30710
rect 4238 30654 4294 30658
rect 4726 32320 4782 32323
rect 4726 32267 4728 32320
rect 4728 32267 4780 32320
rect 4780 32267 4782 32320
rect 4726 32125 4728 32181
rect 4728 32125 4780 32181
rect 4780 32125 4782 32181
rect 4726 31983 4728 32039
rect 4728 31983 4780 32039
rect 4780 31983 4782 32039
rect 4726 31841 4728 31897
rect 4728 31841 4780 31897
rect 4780 31841 4782 31897
rect 4726 31699 4728 31755
rect 4728 31699 4780 31755
rect 4780 31699 4782 31755
rect 4726 31557 4728 31613
rect 4728 31557 4780 31613
rect 4780 31557 4782 31613
rect 4726 31415 4728 31471
rect 4728 31415 4780 31471
rect 4780 31415 4782 31471
rect 4726 31273 4728 31329
rect 4728 31273 4780 31329
rect 4780 31273 4782 31329
rect 4726 31131 4728 31187
rect 4728 31131 4780 31187
rect 4780 31131 4782 31187
rect 4726 30989 4728 31045
rect 4728 30989 4780 31045
rect 4780 30989 4782 31045
rect 4726 30847 4728 30903
rect 4728 30847 4780 30903
rect 4780 30847 4782 30903
rect 4726 30708 4728 30761
rect 4728 30708 4780 30761
rect 4780 30708 4782 30761
rect 4726 30705 4782 30708
rect 5214 32320 5270 32323
rect 5214 32267 5216 32320
rect 5216 32267 5268 32320
rect 5268 32267 5270 32320
rect 5214 32125 5216 32181
rect 5216 32125 5268 32181
rect 5268 32125 5270 32181
rect 5214 31983 5216 32039
rect 5216 31983 5268 32039
rect 5268 31983 5270 32039
rect 5214 31841 5216 31897
rect 5216 31841 5268 31897
rect 5268 31841 5270 31897
rect 5214 31699 5216 31755
rect 5216 31699 5268 31755
rect 5268 31699 5270 31755
rect 5214 31557 5216 31613
rect 5216 31557 5268 31613
rect 5268 31557 5270 31613
rect 5214 31415 5216 31471
rect 5216 31415 5268 31471
rect 5268 31415 5270 31471
rect 5214 31273 5216 31329
rect 5216 31273 5268 31329
rect 5268 31273 5270 31329
rect 5214 31131 5216 31187
rect 5216 31131 5268 31187
rect 5268 31131 5270 31187
rect 5214 30989 5216 31045
rect 5216 30989 5268 31045
rect 5268 30989 5270 31045
rect 5214 30847 5216 30903
rect 5216 30847 5268 30903
rect 5268 30847 5270 30903
rect 5214 30708 5216 30761
rect 5216 30708 5268 30761
rect 5268 30708 5270 30761
rect 5214 30705 5270 30708
rect 5630 32320 5686 32323
rect 5630 32267 5632 32320
rect 5632 32267 5684 32320
rect 5684 32267 5686 32320
rect 5630 32125 5632 32181
rect 5632 32125 5684 32181
rect 5684 32125 5686 32181
rect 5630 31983 5632 32039
rect 5632 31983 5684 32039
rect 5684 31983 5686 32039
rect 5630 31841 5632 31897
rect 5632 31841 5684 31897
rect 5684 31841 5686 31897
rect 5630 31699 5632 31755
rect 5632 31699 5684 31755
rect 5684 31699 5686 31755
rect 5630 31557 5632 31613
rect 5632 31557 5684 31613
rect 5684 31557 5686 31613
rect 5630 31415 5632 31471
rect 5632 31415 5684 31471
rect 5684 31415 5686 31471
rect 5630 31273 5632 31329
rect 5632 31273 5684 31329
rect 5684 31273 5686 31329
rect 5630 31131 5632 31187
rect 5632 31131 5684 31187
rect 5684 31131 5686 31187
rect 5630 30989 5632 31045
rect 5632 30989 5684 31045
rect 5684 30989 5686 31045
rect 5630 30847 5632 30903
rect 5632 30847 5684 30903
rect 5684 30847 5686 30903
rect 5630 30708 5632 30761
rect 5632 30708 5684 30761
rect 5684 30708 5686 30761
rect 5630 30705 5686 30708
rect 7022 32320 7078 32322
rect 7022 32266 7024 32320
rect 7024 32266 7076 32320
rect 7076 32266 7078 32320
rect 7022 32124 7024 32180
rect 7024 32124 7076 32180
rect 7076 32124 7078 32180
rect 7022 31982 7024 32038
rect 7024 31982 7076 32038
rect 7076 31982 7078 32038
rect 7022 31840 7024 31896
rect 7024 31840 7076 31896
rect 7076 31840 7078 31896
rect 7022 31698 7024 31754
rect 7024 31698 7076 31754
rect 7076 31698 7078 31754
rect 7022 31556 7024 31612
rect 7024 31556 7076 31612
rect 7076 31556 7078 31612
rect 7022 31414 7024 31470
rect 7024 31414 7076 31470
rect 7076 31414 7078 31470
rect 7022 31272 7024 31328
rect 7024 31272 7076 31328
rect 7076 31272 7078 31328
rect 7022 31130 7024 31186
rect 7024 31130 7076 31186
rect 7076 31130 7078 31186
rect 7022 30988 7024 31044
rect 7024 30988 7076 31044
rect 7076 30988 7078 31044
rect 7022 30846 7024 30902
rect 7024 30846 7076 30902
rect 7076 30846 7078 30902
rect 7022 30704 7024 30760
rect 7024 30704 7076 30760
rect 7076 30704 7078 30760
rect 2786 30562 2788 30618
rect 2788 30562 2840 30618
rect 2840 30562 2842 30618
rect 7022 30562 7024 30618
rect 7024 30562 7076 30618
rect 7076 30562 7078 30618
rect 2786 30420 2788 30476
rect 2788 30420 2840 30476
rect 2840 30420 2842 30476
rect 2786 30278 2788 30334
rect 2788 30278 2840 30334
rect 2840 30278 2842 30334
rect 2786 30136 2788 30192
rect 2788 30136 2840 30192
rect 2840 30136 2842 30192
rect 175 28141 231 28197
rect 317 28141 373 28197
rect 175 27999 231 28055
rect 317 27999 373 28055
rect 1995 29737 2051 29739
rect 2137 29737 2193 29739
rect 2279 29737 2335 29739
rect 2421 29737 2477 29739
rect 2563 29737 2619 29739
rect 2705 29737 2761 29739
rect 2847 29737 2903 29739
rect 2989 29737 3045 29739
rect 3131 29737 3187 29739
rect 3273 29737 3329 29739
rect 1995 29685 2012 29737
rect 2012 29685 2051 29737
rect 2137 29685 2193 29737
rect 2279 29685 2335 29737
rect 2421 29685 2477 29737
rect 2563 29685 2619 29737
rect 2705 29685 2761 29737
rect 2847 29685 2903 29737
rect 2989 29685 3045 29737
rect 3131 29685 3187 29737
rect 3273 29685 3312 29737
rect 3312 29685 3329 29737
rect 1995 29683 2051 29685
rect 2137 29683 2193 29685
rect 2279 29683 2335 29685
rect 2421 29683 2477 29685
rect 2563 29683 2619 29685
rect 2705 29683 2761 29685
rect 2847 29683 2903 29685
rect 2989 29683 3045 29685
rect 3131 29683 3187 29685
rect 3273 29683 3329 29685
rect 7022 30420 7024 30476
rect 7024 30420 7076 30476
rect 7076 30420 7078 30476
rect 7022 30278 7024 30334
rect 7024 30278 7076 30334
rect 7076 30278 7078 30334
rect 7022 30136 7024 30192
rect 7024 30136 7076 30192
rect 7076 30136 7078 30192
rect 175 27857 231 27913
rect 317 27857 373 27913
rect 175 27715 231 27771
rect 317 27715 373 27771
rect 7997 39944 8053 39946
rect 8139 39944 8195 39946
rect 8281 39944 8337 39946
rect 8423 39944 8479 39946
rect 8565 39944 8621 39946
rect 8707 39944 8763 39946
rect 8849 39944 8905 39946
rect 8991 39944 9047 39946
rect 9133 39944 9189 39946
rect 9275 39944 9331 39946
rect 9417 39944 9473 39946
rect 9559 39944 9615 39946
rect 9701 39944 9757 39946
rect 7997 39892 8053 39944
rect 8139 39892 8195 39944
rect 8281 39892 8337 39944
rect 8423 39892 8479 39944
rect 8565 39892 8621 39944
rect 8707 39892 8763 39944
rect 8849 39892 8905 39944
rect 8991 39892 9047 39944
rect 9133 39892 9189 39944
rect 9275 39892 9331 39944
rect 9417 39892 9473 39944
rect 9559 39892 9615 39944
rect 9701 39892 9720 39944
rect 9720 39892 9757 39944
rect 7997 39890 8053 39892
rect 8139 39890 8195 39892
rect 8281 39890 8337 39892
rect 8423 39890 8479 39892
rect 8565 39890 8621 39892
rect 8707 39890 8763 39892
rect 8849 39890 8905 39892
rect 8991 39890 9047 39892
rect 9133 39890 9189 39892
rect 9275 39890 9331 39892
rect 9417 39890 9473 39892
rect 9559 39890 9615 39892
rect 9701 39890 9757 39892
rect 10337 39358 10339 39414
rect 10339 39358 10391 39414
rect 10391 39358 10393 39414
rect 10337 39216 10339 39272
rect 10339 39216 10391 39272
rect 10391 39216 10393 39272
rect 10337 39074 10339 39130
rect 10339 39074 10391 39130
rect 10391 39074 10393 39130
rect 10337 38932 10339 38988
rect 10339 38932 10391 38988
rect 10391 38932 10393 38988
rect 10337 38790 10339 38846
rect 10339 38790 10391 38846
rect 10391 38790 10393 38846
rect 10337 38648 10339 38704
rect 10339 38648 10391 38704
rect 10391 38648 10393 38704
rect 10337 38506 10339 38562
rect 10339 38506 10391 38562
rect 10391 38506 10393 38562
rect 11210 39358 11212 39414
rect 11212 39358 11264 39414
rect 11264 39358 11266 39414
rect 11210 39216 11212 39272
rect 11212 39216 11264 39272
rect 11264 39216 11266 39272
rect 11210 39074 11212 39130
rect 11212 39074 11264 39130
rect 11264 39074 11266 39130
rect 11210 38932 11212 38988
rect 11212 38932 11264 38988
rect 11264 38932 11266 38988
rect 11210 38790 11212 38846
rect 11212 38790 11264 38846
rect 11264 38790 11266 38846
rect 11210 38648 11212 38704
rect 11212 38648 11264 38704
rect 11264 38648 11266 38704
rect 10337 38364 10393 38420
rect 11210 38506 11212 38562
rect 11212 38506 11264 38562
rect 11264 38506 11266 38562
rect 11210 38364 11266 38420
rect 8681 35576 8737 35612
rect 8681 35556 8735 35576
rect 8735 35556 8737 35576
rect 8681 35414 8737 35470
rect 8681 35272 8737 35328
rect 8681 35130 8737 35186
rect 8681 34988 8737 35044
rect 8681 34846 8737 34902
rect 8681 34704 8737 34760
rect 8681 34562 8737 34618
rect 8681 34420 8737 34476
rect 8681 34278 8737 34334
rect 8681 34136 8737 34192
rect 13191 42542 13247 42598
rect 13303 42542 13359 42598
rect 13415 42542 13471 42598
rect 13191 42430 13247 42486
rect 13303 42430 13359 42486
rect 13415 42430 13471 42486
rect 13191 42318 13247 42374
rect 13303 42318 13359 42374
rect 13415 42318 13471 42374
rect 13191 42206 13247 42262
rect 13303 42206 13359 42262
rect 13415 42206 13471 42262
rect 13191 42094 13247 42150
rect 13303 42094 13359 42150
rect 13415 42094 13471 42150
rect 13191 41982 13247 42038
rect 13303 41982 13359 42038
rect 13415 41982 13471 42038
rect 13191 41870 13247 41926
rect 13303 41870 13359 41926
rect 13415 41870 13471 41926
rect 13191 41758 13247 41814
rect 13303 41758 13359 41814
rect 13415 41758 13471 41814
rect 13191 41646 13247 41702
rect 13303 41646 13359 41702
rect 13415 41646 13471 41702
rect 13191 41534 13247 41590
rect 13303 41534 13359 41590
rect 13415 41534 13471 41590
rect 13191 41422 13247 41478
rect 13303 41422 13359 41478
rect 13415 41422 13471 41478
rect 14410 55341 14466 55397
rect 14552 55341 14608 55397
rect 14694 55341 14750 55397
rect 14410 55199 14466 55255
rect 14552 55199 14608 55255
rect 14694 55199 14750 55255
rect 14410 55057 14466 55113
rect 14552 55057 14608 55113
rect 14694 55057 14750 55113
rect 14410 54915 14466 54971
rect 14552 54915 14608 54971
rect 14694 54915 14750 54971
rect 14410 54773 14466 54829
rect 14552 54773 14608 54829
rect 14694 54773 14750 54829
rect 14410 54631 14466 54687
rect 14552 54631 14608 54687
rect 14694 54631 14750 54687
rect 14410 54489 14466 54545
rect 14552 54489 14608 54545
rect 14694 54489 14750 54545
rect 14410 54347 14466 54403
rect 14552 54347 14608 54403
rect 14694 54347 14750 54403
rect 14410 54205 14466 54261
rect 14552 54205 14608 54261
rect 14694 54205 14750 54261
rect 14410 54063 14466 54119
rect 14552 54063 14608 54119
rect 14694 54063 14750 54119
rect 14952 52180 15008 52197
rect 14952 52141 14954 52180
rect 14954 52141 15006 52180
rect 15006 52141 15008 52180
rect 14952 51999 14954 52055
rect 14954 51999 15006 52055
rect 15006 51999 15008 52055
rect 14952 51857 14954 51913
rect 14954 51857 15006 51913
rect 15006 51857 15008 51913
rect 14952 51715 14954 51771
rect 14954 51715 15006 51771
rect 15006 51715 15008 51771
rect 14952 51573 14954 51629
rect 14954 51573 15006 51629
rect 15006 51573 15008 51629
rect 14952 51431 14954 51487
rect 14954 51431 15006 51487
rect 15006 51431 15008 51487
rect 14952 51289 14954 51345
rect 14954 51289 15006 51345
rect 15006 51289 15008 51345
rect 14952 51147 14954 51203
rect 14954 51147 15006 51203
rect 15006 51147 15008 51203
rect 14952 51005 14954 51061
rect 14954 51005 15006 51061
rect 15006 51005 15008 51061
rect 14952 50880 14954 50919
rect 14954 50880 15006 50919
rect 15006 50880 15008 50919
rect 14952 50863 15008 50880
rect 14410 44141 14466 44197
rect 14552 44141 14608 44197
rect 14694 44141 14750 44197
rect 14410 43999 14466 44055
rect 14552 43999 14608 44055
rect 14694 43999 14750 44055
rect 14410 43857 14466 43913
rect 14552 43857 14608 43913
rect 14694 43857 14750 43913
rect 14410 43715 14466 43771
rect 14552 43715 14608 43771
rect 14694 43715 14750 43771
rect 14410 43573 14466 43629
rect 14552 43573 14608 43629
rect 14694 43573 14750 43629
rect 14410 43431 14466 43487
rect 14552 43431 14608 43487
rect 14694 43431 14750 43487
rect 14410 43289 14466 43345
rect 14552 43289 14608 43345
rect 14694 43289 14750 43345
rect 14410 43147 14466 43203
rect 14552 43147 14608 43203
rect 14694 43147 14750 43203
rect 14410 43005 14466 43061
rect 14552 43005 14608 43061
rect 14694 43005 14750 43061
rect 14410 42863 14466 42919
rect 14552 42863 14608 42919
rect 14694 42863 14750 42919
rect 14410 42541 14466 42597
rect 14552 42541 14608 42597
rect 14694 42541 14750 42597
rect 14410 42399 14466 42455
rect 14552 42399 14608 42455
rect 14694 42399 14750 42455
rect 14410 42257 14466 42313
rect 14552 42257 14608 42313
rect 14694 42257 14750 42313
rect 14410 42115 14466 42171
rect 14552 42115 14608 42171
rect 14694 42115 14750 42171
rect 14410 41973 14466 42029
rect 14552 41973 14608 42029
rect 14694 41973 14750 42029
rect 14410 41831 14466 41887
rect 14552 41831 14608 41887
rect 14694 41831 14750 41887
rect 14410 41689 14466 41745
rect 14552 41689 14608 41745
rect 14694 41689 14750 41745
rect 14410 41547 14466 41603
rect 14552 41547 14608 41603
rect 14694 41547 14750 41603
rect 14410 41405 14466 41461
rect 14552 41405 14608 41461
rect 14694 41405 14750 41461
rect 14410 41263 14466 41319
rect 14552 41263 14608 41319
rect 14694 41263 14750 41319
rect 14410 40941 14466 40997
rect 14552 40941 14608 40997
rect 14694 40941 14750 40997
rect 14410 40799 14466 40855
rect 14552 40799 14608 40855
rect 14694 40799 14750 40855
rect 14410 40657 14466 40713
rect 14552 40657 14608 40713
rect 14694 40657 14750 40713
rect 14410 40515 14466 40571
rect 14552 40515 14608 40571
rect 14694 40515 14750 40571
rect 14410 40373 14466 40429
rect 14552 40373 14608 40429
rect 14694 40373 14750 40429
rect 14410 40231 14466 40287
rect 14552 40231 14608 40287
rect 14694 40231 14750 40287
rect 14410 40089 14466 40145
rect 14552 40089 14608 40145
rect 14694 40089 14750 40145
rect 12758 39944 12814 39946
rect 12900 39944 12956 39946
rect 13042 39944 13098 39946
rect 13184 39944 13240 39946
rect 13326 39944 13382 39946
rect 13468 39944 13524 39946
rect 13610 39944 13666 39946
rect 13752 39944 13808 39946
rect 12758 39892 12784 39944
rect 12784 39892 12814 39944
rect 12900 39892 12956 39944
rect 13042 39892 13098 39944
rect 13184 39892 13240 39944
rect 13326 39892 13382 39944
rect 13468 39892 13524 39944
rect 13610 39892 13666 39944
rect 13752 39892 13772 39944
rect 13772 39892 13808 39944
rect 12758 39890 12814 39892
rect 12900 39890 12956 39892
rect 13042 39890 13098 39892
rect 13184 39890 13240 39892
rect 13326 39890 13382 39892
rect 13468 39890 13524 39892
rect 13610 39890 13666 39892
rect 13752 39890 13808 39892
rect 14410 39947 14466 40003
rect 14552 39947 14608 40003
rect 14694 39947 14750 40003
rect 14410 39805 14466 39861
rect 14552 39805 14608 39861
rect 14694 39805 14750 39861
rect 14410 39663 14466 39719
rect 14552 39663 14608 39719
rect 14694 39663 14750 39719
rect 12416 37741 12472 37797
rect 12558 37741 12614 37797
rect 12416 37599 12472 37655
rect 12558 37599 12614 37655
rect 12416 37457 12472 37513
rect 12558 37457 12614 37513
rect 10435 37198 10491 37200
rect 10577 37198 10633 37200
rect 10719 37198 10775 37200
rect 10861 37198 10917 37200
rect 11003 37198 11059 37200
rect 11145 37198 11201 37200
rect 11287 37198 11343 37200
rect 11429 37198 11485 37200
rect 10435 37146 10491 37198
rect 10577 37146 10633 37198
rect 10719 37146 10775 37198
rect 10861 37146 10917 37198
rect 11003 37146 11059 37198
rect 11145 37146 11201 37198
rect 11287 37146 11343 37198
rect 11429 37146 11485 37198
rect 10435 37144 10491 37146
rect 10577 37144 10633 37146
rect 10719 37144 10775 37146
rect 10861 37144 10917 37146
rect 11003 37144 11059 37146
rect 11145 37144 11201 37146
rect 11287 37144 11343 37146
rect 11429 37144 11485 37146
rect 11008 35660 11064 35716
rect 10110 35576 10166 35612
rect 10110 35556 10112 35576
rect 10112 35556 10164 35576
rect 10164 35556 10166 35576
rect 10110 35414 10112 35470
rect 10112 35414 10164 35470
rect 10164 35414 10166 35470
rect 10110 35272 10112 35328
rect 10112 35272 10164 35328
rect 10164 35272 10166 35328
rect 10110 35130 10112 35186
rect 10112 35130 10164 35186
rect 10164 35130 10166 35186
rect 10110 34988 10112 35044
rect 10112 34988 10164 35044
rect 10164 34988 10166 35044
rect 10110 34846 10112 34902
rect 10112 34846 10164 34902
rect 10164 34846 10166 34902
rect 10110 34704 10112 34760
rect 10112 34704 10164 34760
rect 10164 34704 10166 34760
rect 10110 34562 10112 34618
rect 10112 34562 10164 34618
rect 10164 34562 10166 34618
rect 10110 34420 10112 34476
rect 10112 34420 10164 34476
rect 10164 34420 10166 34476
rect 10110 34278 10112 34334
rect 10112 34278 10164 34334
rect 10164 34278 10166 34334
rect 10110 34172 10112 34192
rect 10112 34172 10164 34192
rect 10164 34172 10166 34192
rect 10110 34136 10166 34172
rect 11008 35518 11010 35574
rect 11010 35518 11062 35574
rect 11062 35518 11064 35574
rect 11008 35376 11010 35432
rect 11010 35376 11062 35432
rect 11062 35376 11064 35432
rect 11008 35234 11010 35290
rect 11010 35234 11062 35290
rect 11062 35234 11064 35290
rect 11008 35092 11010 35148
rect 11010 35092 11062 35148
rect 11062 35092 11064 35148
rect 11008 34950 11010 35006
rect 11010 34950 11062 35006
rect 11062 34950 11064 35006
rect 11008 34808 11010 34864
rect 11010 34808 11062 34864
rect 11062 34808 11064 34864
rect 11008 34666 11010 34722
rect 11010 34666 11062 34722
rect 11062 34666 11064 34722
rect 11008 34524 11010 34580
rect 11010 34524 11062 34580
rect 11062 34524 11064 34580
rect 11008 34382 11010 34438
rect 11010 34382 11062 34438
rect 11062 34382 11064 34438
rect 11008 34240 11010 34296
rect 11010 34240 11062 34296
rect 11062 34240 11064 34296
rect 11008 34098 11010 34154
rect 11010 34098 11062 34154
rect 11062 34098 11064 34154
rect 11008 33956 11010 34012
rect 11010 33956 11062 34012
rect 11062 33956 11064 34012
rect 12416 37315 12472 37371
rect 12558 37315 12614 37371
rect 12416 37173 12472 37229
rect 12558 37173 12614 37229
rect 12416 37031 12472 37087
rect 12558 37031 12614 37087
rect 12416 36889 12472 36945
rect 12558 36889 12614 36945
rect 12416 36747 12472 36803
rect 12558 36747 12614 36803
rect 12416 36605 12472 36661
rect 12558 36605 12614 36661
rect 12416 36463 12472 36519
rect 12558 36463 12614 36519
rect 11906 35576 11962 35612
rect 11906 35556 11908 35576
rect 11908 35556 11960 35576
rect 11960 35556 11962 35576
rect 11906 35414 11908 35470
rect 11908 35414 11960 35470
rect 11960 35414 11962 35470
rect 11906 35272 11908 35328
rect 11908 35272 11960 35328
rect 11960 35272 11962 35328
rect 11906 35130 11908 35186
rect 11908 35130 11960 35186
rect 11960 35130 11962 35186
rect 11906 34988 11908 35044
rect 11908 34988 11960 35044
rect 11960 34988 11962 35044
rect 11906 34846 11908 34902
rect 11908 34846 11960 34902
rect 11960 34846 11962 34902
rect 11906 34704 11908 34760
rect 11908 34704 11960 34760
rect 11960 34704 11962 34760
rect 11906 34562 11908 34618
rect 11908 34562 11960 34618
rect 11960 34562 11962 34618
rect 11906 34420 11908 34476
rect 11908 34420 11960 34476
rect 11960 34420 11962 34476
rect 11906 34278 11908 34334
rect 11908 34278 11960 34334
rect 11960 34278 11962 34334
rect 11906 34172 11908 34192
rect 11908 34172 11960 34192
rect 11960 34172 11962 34192
rect 11906 34136 11962 34172
rect 11008 33814 11010 33870
rect 11010 33814 11062 33870
rect 11062 33814 11064 33870
rect 11008 33672 11010 33728
rect 11010 33672 11062 33728
rect 11062 33672 11064 33728
rect 11008 33530 11010 33586
rect 11010 33530 11062 33586
rect 11062 33530 11064 33586
rect 11008 33388 11010 33444
rect 11010 33388 11062 33444
rect 11062 33388 11064 33444
rect 11008 33246 11010 33302
rect 11010 33246 11062 33302
rect 11062 33246 11064 33302
rect 11008 32479 11064 32535
rect 14952 37780 15008 37797
rect 14952 37741 14954 37780
rect 14954 37741 15006 37780
rect 15006 37741 15008 37780
rect 14952 37599 14954 37655
rect 14954 37599 15006 37655
rect 15006 37599 15008 37655
rect 14952 37457 14954 37513
rect 14954 37457 15006 37513
rect 15006 37457 15008 37513
rect 14952 37315 14954 37371
rect 14954 37315 15006 37371
rect 15006 37315 15008 37371
rect 14952 37173 14954 37229
rect 14954 37173 15006 37229
rect 15006 37173 15008 37229
rect 14952 37031 14954 37087
rect 14954 37031 15006 37087
rect 15006 37031 15008 37087
rect 14952 36889 14954 36945
rect 14954 36889 15006 36945
rect 15006 36889 15008 36945
rect 14952 36747 14954 36803
rect 14954 36747 15006 36803
rect 15006 36747 15008 36803
rect 14952 36605 14954 36661
rect 14954 36605 15006 36661
rect 15006 36605 15008 36661
rect 14952 36480 14954 36519
rect 14954 36480 15006 36519
rect 15006 36480 15008 36519
rect 14952 36463 15008 36480
rect 14410 32922 14466 32978
rect 14552 32922 14566 32978
rect 14566 32922 14608 32978
rect 14694 32922 14750 32978
rect 14410 32780 14466 32836
rect 14552 32780 14566 32836
rect 14566 32780 14608 32836
rect 14694 32780 14750 32836
rect 14410 32638 14466 32694
rect 14552 32638 14566 32694
rect 14566 32638 14608 32694
rect 14694 32638 14750 32694
rect 11008 32337 11010 32393
rect 11010 32337 11062 32393
rect 11062 32337 11064 32393
rect 7986 32320 8042 32322
rect 7986 32266 7988 32320
rect 7988 32266 8040 32320
rect 8040 32266 8042 32320
rect 7986 32124 7988 32180
rect 7988 32124 8040 32180
rect 8040 32124 8042 32180
rect 7986 31982 7988 32038
rect 7988 31982 8040 32038
rect 8040 31982 8042 32038
rect 7986 31840 7988 31896
rect 7988 31840 8040 31896
rect 8040 31840 8042 31896
rect 7986 31698 7988 31754
rect 7988 31698 8040 31754
rect 8040 31698 8042 31754
rect 7986 31556 7988 31612
rect 7988 31556 8040 31612
rect 8040 31556 8042 31612
rect 7986 31414 7988 31470
rect 7988 31414 8040 31470
rect 8040 31414 8042 31470
rect 7986 31272 7988 31328
rect 7988 31272 8040 31328
rect 8040 31272 8042 31328
rect 7986 31130 7988 31186
rect 7988 31130 8040 31186
rect 8040 31130 8042 31186
rect 7986 30988 7988 31044
rect 7988 30988 8040 31044
rect 8040 30988 8042 31044
rect 7986 30846 7988 30902
rect 7988 30846 8040 30902
rect 8040 30846 8042 30902
rect 7986 30704 7988 30760
rect 7988 30704 8040 30760
rect 8040 30704 8042 30760
rect 9378 32320 9434 32323
rect 9378 32267 9380 32320
rect 9380 32267 9432 32320
rect 9432 32267 9434 32320
rect 9378 32125 9380 32181
rect 9380 32125 9432 32181
rect 9432 32125 9434 32181
rect 9378 31983 9380 32039
rect 9380 31983 9432 32039
rect 9432 31983 9434 32039
rect 9378 31841 9380 31897
rect 9380 31841 9432 31897
rect 9432 31841 9434 31897
rect 9378 31699 9380 31755
rect 9380 31699 9432 31755
rect 9432 31699 9434 31755
rect 9378 31557 9380 31613
rect 9380 31557 9432 31613
rect 9432 31557 9434 31613
rect 9378 31415 9380 31471
rect 9380 31415 9432 31471
rect 9432 31415 9434 31471
rect 9378 31273 9380 31329
rect 9380 31273 9432 31329
rect 9432 31273 9434 31329
rect 9378 31131 9380 31187
rect 9380 31131 9432 31187
rect 9432 31131 9434 31187
rect 9378 30989 9380 31045
rect 9380 30989 9432 31045
rect 9432 30989 9434 31045
rect 9378 30847 9380 30903
rect 9380 30847 9432 30903
rect 9432 30847 9434 30903
rect 9378 30708 9380 30761
rect 9380 30708 9432 30761
rect 9432 30708 9434 30761
rect 9378 30705 9434 30708
rect 9794 32320 9850 32323
rect 9794 32267 9796 32320
rect 9796 32267 9848 32320
rect 9848 32267 9850 32320
rect 9794 32125 9796 32181
rect 9796 32125 9848 32181
rect 9848 32125 9850 32181
rect 9794 31983 9796 32039
rect 9796 31983 9848 32039
rect 9848 31983 9850 32039
rect 9794 31841 9796 31897
rect 9796 31841 9848 31897
rect 9848 31841 9850 31897
rect 9794 31699 9796 31755
rect 9796 31699 9848 31755
rect 9848 31699 9850 31755
rect 9794 31557 9796 31613
rect 9796 31557 9848 31613
rect 9848 31557 9850 31613
rect 9794 31415 9796 31471
rect 9796 31415 9848 31471
rect 9848 31415 9850 31471
rect 9794 31273 9796 31329
rect 9796 31273 9848 31329
rect 9848 31273 9850 31329
rect 9794 31131 9796 31187
rect 9796 31131 9848 31187
rect 9848 31131 9850 31187
rect 9794 30989 9796 31045
rect 9796 30989 9848 31045
rect 9848 30989 9850 31045
rect 9794 30847 9796 30903
rect 9796 30847 9848 30903
rect 9848 30847 9850 30903
rect 9794 30708 9796 30761
rect 9796 30708 9848 30761
rect 9848 30708 9850 30761
rect 9794 30705 9850 30708
rect 10282 32320 10338 32323
rect 10282 32267 10284 32320
rect 10284 32267 10336 32320
rect 10336 32267 10338 32320
rect 10282 32125 10284 32181
rect 10284 32125 10336 32181
rect 10336 32125 10338 32181
rect 10282 31983 10284 32039
rect 10284 31983 10336 32039
rect 10336 31983 10338 32039
rect 10282 31841 10284 31897
rect 10284 31841 10336 31897
rect 10336 31841 10338 31897
rect 10282 31699 10284 31755
rect 10284 31699 10336 31755
rect 10336 31699 10338 31755
rect 10282 31557 10284 31613
rect 10284 31557 10336 31613
rect 10336 31557 10338 31613
rect 10282 31415 10284 31471
rect 10284 31415 10336 31471
rect 10336 31415 10338 31471
rect 10282 31273 10284 31329
rect 10284 31273 10336 31329
rect 10336 31273 10338 31329
rect 10282 31131 10284 31187
rect 10284 31131 10336 31187
rect 10336 31131 10338 31187
rect 10282 30989 10284 31045
rect 10284 30989 10336 31045
rect 10336 30989 10338 31045
rect 10282 30847 10284 30903
rect 10284 30847 10336 30903
rect 10336 30847 10338 30903
rect 10282 30708 10284 30761
rect 10284 30708 10336 30761
rect 10336 30708 10338 30761
rect 10282 30705 10338 30708
rect 10770 32270 10826 32272
rect 10770 32216 10772 32270
rect 10772 32216 10824 32270
rect 10824 32216 10826 32270
rect 10770 32074 10772 32130
rect 10772 32074 10824 32130
rect 10824 32074 10826 32130
rect 10770 31932 10772 31988
rect 10772 31932 10824 31988
rect 10824 31932 10826 31988
rect 10770 31790 10772 31846
rect 10772 31790 10824 31846
rect 10824 31790 10826 31846
rect 10770 31648 10772 31704
rect 10772 31648 10824 31704
rect 10824 31648 10826 31704
rect 10770 31506 10772 31562
rect 10772 31506 10824 31562
rect 10824 31506 10826 31562
rect 10770 31364 10772 31420
rect 10772 31364 10824 31420
rect 10824 31364 10826 31420
rect 10770 31222 10772 31278
rect 10772 31222 10824 31278
rect 10824 31222 10826 31278
rect 10770 31080 10772 31136
rect 10772 31080 10824 31136
rect 10824 31080 10826 31136
rect 10770 30938 10772 30994
rect 10772 30938 10824 30994
rect 10824 30938 10826 30994
rect 10770 30796 10772 30852
rect 10772 30796 10824 30852
rect 10824 30796 10826 30852
rect 10770 30658 10772 30710
rect 10772 30658 10824 30710
rect 10824 30658 10826 30710
rect 10770 30654 10826 30658
rect 14410 32496 14466 32552
rect 14552 32496 14566 32552
rect 14566 32496 14608 32552
rect 14694 32496 14750 32552
rect 14410 32354 14466 32410
rect 14552 32354 14566 32410
rect 14566 32354 14608 32410
rect 14694 32354 14750 32410
rect 11008 32195 11010 32251
rect 11010 32195 11062 32251
rect 11062 32195 11064 32251
rect 11008 32053 11010 32109
rect 11010 32053 11062 32109
rect 11062 32053 11064 32109
rect 11008 31911 11010 31967
rect 11010 31911 11062 31967
rect 11062 31911 11064 31967
rect 11008 31769 11010 31825
rect 11010 31769 11062 31825
rect 11062 31769 11064 31825
rect 11008 31627 11010 31683
rect 11010 31627 11062 31683
rect 11062 31627 11064 31683
rect 11008 31485 11010 31541
rect 11010 31485 11062 31541
rect 11062 31485 11064 31541
rect 11008 31343 11010 31399
rect 11010 31343 11062 31399
rect 11062 31343 11064 31399
rect 11008 31201 11010 31257
rect 11010 31201 11062 31257
rect 11062 31201 11064 31257
rect 11008 31059 11010 31115
rect 11010 31059 11062 31115
rect 11062 31059 11064 31115
rect 11008 30917 11010 30973
rect 11010 30917 11062 30973
rect 11062 30917 11064 30973
rect 11008 30775 11010 30831
rect 11010 30775 11062 30831
rect 11062 30775 11064 30831
rect 11008 30635 11010 30689
rect 11010 30635 11062 30689
rect 11062 30635 11064 30689
rect 11008 30633 11064 30635
rect 11246 32270 11302 32272
rect 11246 32216 11248 32270
rect 11248 32216 11300 32270
rect 11300 32216 11302 32270
rect 11246 32074 11248 32130
rect 11248 32074 11300 32130
rect 11300 32074 11302 32130
rect 11246 31932 11248 31988
rect 11248 31932 11300 31988
rect 11300 31932 11302 31988
rect 11246 31790 11248 31846
rect 11248 31790 11300 31846
rect 11300 31790 11302 31846
rect 11246 31648 11248 31704
rect 11248 31648 11300 31704
rect 11300 31648 11302 31704
rect 11246 31506 11248 31562
rect 11248 31506 11300 31562
rect 11300 31506 11302 31562
rect 11246 31364 11248 31420
rect 11248 31364 11300 31420
rect 11300 31364 11302 31420
rect 11246 31222 11248 31278
rect 11248 31222 11300 31278
rect 11300 31222 11302 31278
rect 11246 31080 11248 31136
rect 11248 31080 11300 31136
rect 11300 31080 11302 31136
rect 11246 30938 11248 30994
rect 11248 30938 11300 30994
rect 11300 30938 11302 30994
rect 11246 30796 11248 30852
rect 11248 30796 11300 30852
rect 11300 30796 11302 30852
rect 11246 30658 11248 30710
rect 11248 30658 11300 30710
rect 11300 30658 11302 30710
rect 11246 30654 11302 30658
rect 11734 32320 11790 32323
rect 11734 32267 11736 32320
rect 11736 32267 11788 32320
rect 11788 32267 11790 32320
rect 11734 32125 11736 32181
rect 11736 32125 11788 32181
rect 11788 32125 11790 32181
rect 11734 31983 11736 32039
rect 11736 31983 11788 32039
rect 11788 31983 11790 32039
rect 11734 31841 11736 31897
rect 11736 31841 11788 31897
rect 11788 31841 11790 31897
rect 11734 31699 11736 31755
rect 11736 31699 11788 31755
rect 11788 31699 11790 31755
rect 11734 31557 11736 31613
rect 11736 31557 11788 31613
rect 11788 31557 11790 31613
rect 11734 31415 11736 31471
rect 11736 31415 11788 31471
rect 11788 31415 11790 31471
rect 11734 31273 11736 31329
rect 11736 31273 11788 31329
rect 11788 31273 11790 31329
rect 11734 31131 11736 31187
rect 11736 31131 11788 31187
rect 11788 31131 11790 31187
rect 11734 30989 11736 31045
rect 11736 30989 11788 31045
rect 11788 30989 11790 31045
rect 11734 30847 11736 30903
rect 11736 30847 11788 30903
rect 11788 30847 11790 30903
rect 11734 30708 11736 30761
rect 11736 30708 11788 30761
rect 11788 30708 11790 30761
rect 11734 30705 11790 30708
rect 12222 32320 12278 32322
rect 12222 32266 12224 32320
rect 12224 32266 12276 32320
rect 12276 32266 12278 32320
rect 12222 32124 12224 32180
rect 12224 32124 12276 32180
rect 12276 32124 12278 32180
rect 12222 31982 12224 32038
rect 12224 31982 12276 32038
rect 12276 31982 12278 32038
rect 12222 31840 12224 31896
rect 12224 31840 12276 31896
rect 12276 31840 12278 31896
rect 12222 31698 12224 31754
rect 12224 31698 12276 31754
rect 12276 31698 12278 31754
rect 12222 31556 12224 31612
rect 12224 31556 12276 31612
rect 12276 31556 12278 31612
rect 12222 31414 12224 31470
rect 12224 31414 12276 31470
rect 12276 31414 12278 31470
rect 12222 31272 12224 31328
rect 12224 31272 12276 31328
rect 12276 31272 12278 31328
rect 12222 31130 12224 31186
rect 12224 31130 12276 31186
rect 12276 31130 12278 31186
rect 12222 30988 12224 31044
rect 12224 30988 12276 31044
rect 12276 30988 12278 31044
rect 12222 30846 12224 30902
rect 12224 30846 12276 30902
rect 12276 30846 12278 30902
rect 12222 30704 12224 30760
rect 12224 30704 12276 30760
rect 12276 30704 12278 30760
rect 7986 30562 7988 30618
rect 7988 30562 8040 30618
rect 8040 30562 8042 30618
rect 12222 30562 12224 30618
rect 12224 30562 12276 30618
rect 12276 30562 12278 30618
rect 7986 30420 7988 30476
rect 7988 30420 8040 30476
rect 8040 30420 8042 30476
rect 7986 30278 7988 30334
rect 7988 30278 8040 30334
rect 8040 30278 8042 30334
rect 7986 30136 7988 30192
rect 7988 30136 8040 30192
rect 8040 30136 8042 30192
rect 12222 30420 12224 30476
rect 12224 30420 12276 30476
rect 12276 30420 12278 30476
rect 12222 30278 12224 30334
rect 12224 30278 12276 30334
rect 12276 30278 12278 30334
rect 12222 30136 12224 30192
rect 12224 30136 12276 30192
rect 12276 30136 12278 30192
rect 12638 32320 12694 32322
rect 12638 32266 12640 32320
rect 12640 32266 12692 32320
rect 12692 32266 12694 32320
rect 12638 32124 12640 32180
rect 12640 32124 12692 32180
rect 12692 32124 12694 32180
rect 12638 31982 12640 32038
rect 12640 31982 12692 32038
rect 12692 31982 12694 32038
rect 12638 31840 12640 31896
rect 12640 31840 12692 31896
rect 12692 31840 12694 31896
rect 12638 31698 12640 31754
rect 12640 31698 12692 31754
rect 12692 31698 12694 31754
rect 12638 31556 12640 31612
rect 12640 31556 12692 31612
rect 12692 31556 12694 31612
rect 12638 31414 12640 31470
rect 12640 31414 12692 31470
rect 12692 31414 12694 31470
rect 12638 31272 12640 31328
rect 12640 31272 12692 31328
rect 12692 31272 12694 31328
rect 12638 31130 12640 31186
rect 12640 31130 12692 31186
rect 12692 31130 12694 31186
rect 12638 30988 12640 31044
rect 12640 30988 12692 31044
rect 12692 30988 12694 31044
rect 12638 30846 12640 30902
rect 12640 30846 12692 30902
rect 12692 30846 12694 30902
rect 12638 30704 12640 30760
rect 12640 30704 12692 30760
rect 12692 30704 12694 30760
rect 12638 30562 12640 30618
rect 12640 30562 12692 30618
rect 12692 30562 12694 30618
rect 12638 30420 12640 30476
rect 12640 30420 12692 30476
rect 12692 30420 12694 30476
rect 12638 30278 12640 30334
rect 12640 30278 12692 30334
rect 12692 30278 12694 30334
rect 14030 32320 14086 32322
rect 14030 32266 14032 32320
rect 14032 32266 14084 32320
rect 14084 32266 14086 32320
rect 14030 32124 14032 32180
rect 14032 32124 14084 32180
rect 14084 32124 14086 32180
rect 14030 31982 14032 32038
rect 14032 31982 14084 32038
rect 14084 31982 14086 32038
rect 14030 31840 14032 31896
rect 14032 31840 14084 31896
rect 14084 31840 14086 31896
rect 14030 31698 14032 31754
rect 14032 31698 14084 31754
rect 14084 31698 14086 31754
rect 14030 31556 14032 31612
rect 14032 31556 14084 31612
rect 14084 31556 14086 31612
rect 14030 31414 14032 31470
rect 14032 31414 14084 31470
rect 14084 31414 14086 31470
rect 14030 31272 14032 31328
rect 14032 31272 14084 31328
rect 14084 31272 14086 31328
rect 14030 31130 14032 31186
rect 14032 31130 14084 31186
rect 14084 31130 14086 31186
rect 14030 30988 14032 31044
rect 14032 30988 14084 31044
rect 14084 30988 14086 31044
rect 14030 30846 14032 30902
rect 14032 30846 14084 30902
rect 14084 30846 14086 30902
rect 14030 30704 14032 30760
rect 14032 30704 14084 30760
rect 14084 30704 14086 30760
rect 14030 30562 14032 30618
rect 14032 30562 14084 30618
rect 14084 30562 14086 30618
rect 14030 30420 14032 30476
rect 14032 30420 14084 30476
rect 14084 30420 14086 30476
rect 12638 30136 12640 30192
rect 12640 30136 12692 30192
rect 12692 30136 12694 30192
rect 11932 29737 11988 29739
rect 12074 29737 12130 29739
rect 12216 29737 12272 29739
rect 12358 29737 12414 29739
rect 12500 29737 12556 29739
rect 12642 29737 12698 29739
rect 12784 29737 12840 29739
rect 12926 29737 12982 29739
rect 13068 29737 13124 29739
rect 13210 29737 13266 29739
rect 11932 29685 11949 29737
rect 11949 29685 11988 29737
rect 12074 29685 12130 29737
rect 12216 29685 12272 29737
rect 12358 29685 12414 29737
rect 12500 29685 12556 29737
rect 12642 29685 12698 29737
rect 12784 29685 12840 29737
rect 12926 29685 12982 29737
rect 13068 29685 13124 29737
rect 13210 29685 13249 29737
rect 13249 29685 13266 29737
rect 11932 29683 11988 29685
rect 12074 29683 12130 29685
rect 12216 29683 12272 29685
rect 12358 29683 12414 29685
rect 12500 29683 12556 29685
rect 12642 29683 12698 29685
rect 12784 29683 12840 29685
rect 12926 29683 12982 29685
rect 13068 29683 13124 29685
rect 13210 29683 13266 29685
rect 14030 30278 14032 30334
rect 14032 30278 14084 30334
rect 14084 30278 14086 30334
rect 14030 30136 14032 30192
rect 14032 30136 14084 30192
rect 14084 30136 14086 30192
rect 14410 32212 14466 32268
rect 14552 32212 14566 32268
rect 14566 32212 14608 32268
rect 14694 32212 14750 32268
rect 14410 32070 14466 32126
rect 14552 32070 14566 32126
rect 14566 32070 14608 32126
rect 14694 32070 14750 32126
rect 14410 31928 14466 31984
rect 14552 31928 14566 31984
rect 14566 31928 14608 31984
rect 14694 31928 14750 31984
rect 14410 31786 14466 31842
rect 14552 31786 14566 31842
rect 14566 31786 14608 31842
rect 14694 31786 14750 31842
rect 14410 31644 14466 31700
rect 14552 31644 14566 31700
rect 14566 31644 14608 31700
rect 14694 31644 14750 31700
rect 14410 31502 14466 31558
rect 14552 31502 14566 31558
rect 14566 31502 14608 31558
rect 14694 31502 14750 31558
rect 14410 31360 14466 31416
rect 14552 31360 14566 31416
rect 14566 31360 14608 31416
rect 14694 31360 14750 31416
rect 14410 31218 14466 31274
rect 14552 31218 14566 31274
rect 14566 31218 14608 31274
rect 14694 31218 14750 31274
rect 14410 31076 14466 31132
rect 14552 31076 14566 31132
rect 14566 31076 14608 31132
rect 14694 31076 14750 31132
rect 14410 30934 14466 30990
rect 14552 30934 14566 30990
rect 14566 30934 14608 30990
rect 14694 30934 14750 30990
rect 14410 30792 14466 30848
rect 14552 30792 14566 30848
rect 14566 30792 14608 30848
rect 14694 30792 14750 30848
rect 14410 30650 14466 30706
rect 14552 30650 14566 30706
rect 14566 30650 14608 30706
rect 14694 30650 14750 30706
rect 14410 30508 14466 30564
rect 14552 30508 14566 30564
rect 14566 30508 14608 30564
rect 14694 30508 14750 30564
rect 14410 30366 14466 30422
rect 14552 30366 14566 30422
rect 14566 30366 14608 30422
rect 14694 30366 14750 30422
rect 14410 30224 14466 30280
rect 14552 30224 14566 30280
rect 14566 30224 14608 30280
rect 14694 30224 14750 30280
rect 14410 30082 14466 30138
rect 14552 30082 14566 30138
rect 14566 30082 14608 30138
rect 14694 30082 14750 30138
rect 14410 29741 14466 29797
rect 14552 29741 14566 29797
rect 14566 29741 14608 29797
rect 14694 29741 14750 29797
rect 14410 29599 14466 29655
rect 14552 29599 14608 29655
rect 14694 29599 14750 29655
rect 14410 29457 14466 29513
rect 14552 29457 14608 29513
rect 14694 29457 14750 29513
rect 14410 29315 14466 29371
rect 14552 29315 14608 29371
rect 14694 29315 14750 29371
rect 14410 29173 14466 29229
rect 14552 29173 14608 29229
rect 14694 29173 14750 29229
rect 14410 29031 14466 29087
rect 14552 29031 14608 29087
rect 14694 29031 14750 29087
rect 14410 28889 14466 28945
rect 14552 28889 14608 28945
rect 14694 28889 14750 28945
rect 14410 28747 14466 28803
rect 14552 28747 14608 28803
rect 14694 28747 14750 28803
rect 14410 28605 14466 28661
rect 14552 28605 14608 28661
rect 14694 28605 14750 28661
rect 14410 28463 14466 28519
rect 14552 28463 14608 28519
rect 14694 28463 14750 28519
rect 175 27573 231 27629
rect 317 27573 373 27629
rect 175 27431 231 27487
rect 317 27431 373 27487
rect 175 27289 231 27345
rect 317 27289 373 27345
rect 175 27147 231 27203
rect 317 27147 373 27203
rect 175 27005 231 27061
rect 317 27005 373 27061
rect 175 26863 231 26919
rect 317 26863 373 26919
rect 14410 26522 14466 26578
rect 14552 26522 14608 26578
rect 14694 26522 14750 26578
rect 14410 26380 14466 26436
rect 14552 26380 14608 26436
rect 14694 26380 14750 26436
rect 14410 26238 14466 26294
rect 14552 26238 14608 26294
rect 14694 26238 14750 26294
rect 14410 26096 14466 26152
rect 14552 26096 14608 26152
rect 14694 26096 14750 26152
rect 14410 25954 14466 26010
rect 14552 25954 14608 26010
rect 14694 25954 14750 26010
rect 14410 25812 14466 25868
rect 14552 25812 14608 25868
rect 14694 25812 14750 25868
rect 14410 25670 14466 25726
rect 14552 25670 14608 25726
rect 14694 25670 14750 25726
rect 14410 25528 14466 25584
rect 14552 25528 14608 25584
rect 14694 25528 14750 25584
rect 14410 25386 14466 25442
rect 14552 25386 14608 25442
rect 14694 25386 14750 25442
rect 14410 25244 14466 25300
rect 14552 25244 14608 25300
rect 14694 25244 14750 25300
rect 14410 25102 14466 25158
rect 14552 25102 14608 25158
rect 14694 25102 14750 25158
rect 14410 24960 14466 25016
rect 14552 24960 14608 25016
rect 14694 24960 14750 25016
rect 14410 24818 14466 24874
rect 14552 24818 14608 24874
rect 14694 24818 14750 24874
rect 14410 24676 14466 24732
rect 14552 24676 14608 24732
rect 14694 24676 14750 24732
rect 14410 24534 14466 24590
rect 14552 24534 14608 24590
rect 14694 24534 14750 24590
rect 14410 24392 14466 24448
rect 14552 24392 14608 24448
rect 14694 24392 14750 24448
rect 14410 24250 14466 24306
rect 14552 24250 14608 24306
rect 14694 24250 14750 24306
rect 14410 24108 14466 24164
rect 14552 24108 14608 24164
rect 14694 24108 14750 24164
rect 14410 23966 14466 24022
rect 14552 23966 14608 24022
rect 14694 23966 14750 24022
rect 14410 23824 14466 23880
rect 14552 23824 14608 23880
rect 14694 23824 14750 23880
rect 14410 23682 14466 23738
rect 14552 23682 14608 23738
rect 14694 23682 14750 23738
rect 14410 23322 14466 23378
rect 14552 23322 14608 23378
rect 14694 23322 14750 23378
rect 14410 23180 14466 23236
rect 14552 23180 14608 23236
rect 14694 23180 14750 23236
rect 14410 23038 14466 23094
rect 14552 23038 14608 23094
rect 14694 23038 14750 23094
rect 14410 22896 14466 22952
rect 14552 22896 14608 22952
rect 14694 22896 14750 22952
rect 14410 22754 14466 22810
rect 14552 22754 14608 22810
rect 14694 22754 14750 22810
rect 14410 22612 14466 22668
rect 14552 22612 14608 22668
rect 14694 22612 14750 22668
rect 14410 22470 14466 22526
rect 14552 22470 14608 22526
rect 14694 22470 14750 22526
rect 14410 22328 14466 22384
rect 14552 22328 14608 22384
rect 14694 22328 14750 22384
rect 14410 22186 14466 22242
rect 14552 22186 14608 22242
rect 14694 22186 14750 22242
rect 14410 22044 14466 22100
rect 14552 22044 14608 22100
rect 14694 22044 14750 22100
rect 14410 21902 14466 21958
rect 14552 21902 14608 21958
rect 14694 21902 14750 21958
rect 14410 21760 14466 21816
rect 14552 21760 14608 21816
rect 14694 21760 14750 21816
rect 14410 21618 14466 21674
rect 14552 21618 14608 21674
rect 14694 21618 14750 21674
rect 14410 21476 14466 21532
rect 14552 21476 14608 21532
rect 14694 21476 14750 21532
rect 14410 21334 14466 21390
rect 14552 21334 14608 21390
rect 14694 21334 14750 21390
rect 14410 21192 14466 21248
rect 14552 21192 14608 21248
rect 14694 21192 14750 21248
rect 14410 21050 14466 21106
rect 14552 21050 14608 21106
rect 14694 21050 14750 21106
rect 14410 20908 14466 20964
rect 14552 20908 14608 20964
rect 14694 20908 14750 20964
rect 14410 20766 14466 20822
rect 14552 20766 14608 20822
rect 14694 20766 14750 20822
rect 14410 20624 14466 20680
rect 14552 20624 14608 20680
rect 14694 20624 14750 20680
rect 14410 20482 14466 20538
rect 14552 20482 14608 20538
rect 14694 20482 14750 20538
rect 14410 20122 14466 20178
rect 14552 20122 14608 20178
rect 14694 20122 14750 20178
rect 14410 19980 14466 20036
rect 14552 19980 14608 20036
rect 14694 19980 14750 20036
rect 14410 19838 14466 19894
rect 14552 19838 14608 19894
rect 14694 19838 14750 19894
rect 14410 19696 14466 19752
rect 14552 19696 14608 19752
rect 14694 19696 14750 19752
rect 14410 19554 14466 19610
rect 14552 19554 14608 19610
rect 14694 19554 14750 19610
rect 14410 19412 14466 19468
rect 14552 19412 14608 19468
rect 14694 19412 14750 19468
rect 14410 19270 14466 19326
rect 14552 19270 14608 19326
rect 14694 19270 14750 19326
rect 14410 19128 14466 19184
rect 14552 19128 14608 19184
rect 14694 19128 14750 19184
rect 14410 18986 14466 19042
rect 14552 18986 14608 19042
rect 14694 18986 14750 19042
rect 14410 18844 14466 18900
rect 14552 18844 14608 18900
rect 14694 18844 14750 18900
rect 14410 18702 14466 18758
rect 14552 18702 14608 18758
rect 14694 18702 14750 18758
rect 14410 18560 14466 18616
rect 14552 18560 14608 18616
rect 14694 18560 14750 18616
rect 14410 18418 14466 18474
rect 14552 18418 14608 18474
rect 14694 18418 14750 18474
rect 14410 18276 14466 18332
rect 14552 18276 14608 18332
rect 14694 18276 14750 18332
rect 14410 18134 14466 18190
rect 14552 18134 14608 18190
rect 14694 18134 14750 18190
rect 14410 17992 14466 18048
rect 14552 17992 14608 18048
rect 14694 17992 14750 18048
rect 14410 17850 14466 17906
rect 14552 17850 14608 17906
rect 14694 17850 14750 17906
rect 14410 17708 14466 17764
rect 14552 17708 14608 17764
rect 14694 17708 14750 17764
rect 14410 17566 14466 17622
rect 14552 17566 14608 17622
rect 14694 17566 14750 17622
rect 14410 17424 14466 17480
rect 14552 17424 14608 17480
rect 14694 17424 14750 17480
rect 14410 17282 14466 17338
rect 14552 17282 14608 17338
rect 14694 17282 14750 17338
rect 14410 16922 14466 16978
rect 14552 16922 14608 16978
rect 14694 16922 14750 16978
rect 14410 16780 14466 16836
rect 14552 16780 14608 16836
rect 14694 16780 14750 16836
rect 14410 16638 14466 16694
rect 14552 16638 14608 16694
rect 14694 16638 14750 16694
rect 14410 16496 14466 16552
rect 14552 16496 14608 16552
rect 14694 16496 14750 16552
rect 14410 16354 14466 16410
rect 14552 16354 14608 16410
rect 14694 16354 14750 16410
rect 14410 16212 14466 16268
rect 14552 16212 14608 16268
rect 14694 16212 14750 16268
rect 14410 16070 14466 16126
rect 14552 16070 14608 16126
rect 14694 16070 14750 16126
rect 14410 15928 14466 15984
rect 14552 15928 14608 15984
rect 14694 15928 14750 15984
rect 14410 15786 14466 15842
rect 14552 15786 14608 15842
rect 14694 15786 14750 15842
rect 14410 15644 14466 15700
rect 14552 15644 14608 15700
rect 14694 15644 14750 15700
rect 14410 15502 14466 15558
rect 14552 15502 14608 15558
rect 14694 15502 14750 15558
rect 14410 15360 14466 15416
rect 14552 15360 14608 15416
rect 14694 15360 14750 15416
rect 14410 15218 14466 15274
rect 14552 15218 14608 15274
rect 14694 15218 14750 15274
rect 14410 15076 14466 15132
rect 14552 15076 14608 15132
rect 14694 15076 14750 15132
rect 14410 14934 14466 14990
rect 14552 14934 14608 14990
rect 14694 14934 14750 14990
rect 14410 14792 14466 14848
rect 14552 14792 14608 14848
rect 14694 14792 14750 14848
rect 14410 14650 14466 14706
rect 14552 14650 14608 14706
rect 14694 14650 14750 14706
rect 14410 14508 14466 14564
rect 14552 14508 14608 14564
rect 14694 14508 14750 14564
rect 14410 14366 14466 14422
rect 14552 14366 14608 14422
rect 14694 14366 14750 14422
rect 14410 14224 14466 14280
rect 14552 14224 14608 14280
rect 14694 14224 14750 14280
rect 14410 14082 14466 14138
rect 14552 14082 14608 14138
rect 14694 14082 14750 14138
rect 175 10522 231 10578
rect 317 10522 373 10578
rect 175 10380 231 10436
rect 317 10380 373 10436
rect 175 10238 231 10294
rect 317 10238 373 10294
rect 175 10096 231 10152
rect 317 10096 373 10152
rect 175 9954 231 10010
rect 317 9954 373 10010
rect 175 9812 231 9868
rect 317 9812 373 9868
rect 175 9670 231 9726
rect 317 9670 373 9726
rect 175 9528 231 9584
rect 317 9528 373 9584
rect 175 9386 231 9442
rect 317 9386 373 9442
rect 175 9244 231 9300
rect 317 9244 373 9300
rect 175 9102 231 9158
rect 317 9102 373 9158
rect 175 8960 231 9016
rect 317 8960 373 9016
rect 175 8818 231 8874
rect 317 8818 373 8874
rect 175 8676 231 8732
rect 317 8676 373 8732
rect 175 8534 231 8590
rect 317 8534 373 8590
rect 175 8392 231 8448
rect 317 8392 373 8448
rect 175 8250 231 8306
rect 317 8250 373 8306
rect 175 8108 231 8164
rect 317 8108 373 8164
rect 175 7966 231 8022
rect 317 7966 373 8022
rect 175 7824 231 7880
rect 317 7824 373 7880
rect 175 7682 231 7738
rect 317 7682 373 7738
rect 175 7322 231 7378
rect 317 7322 373 7378
rect 175 7180 231 7236
rect 317 7180 373 7236
rect 175 7038 231 7094
rect 317 7038 373 7094
rect 175 6896 231 6952
rect 317 6896 373 6952
rect 175 6754 231 6810
rect 317 6754 373 6810
rect 175 6612 231 6668
rect 317 6612 373 6668
rect 175 6470 231 6526
rect 317 6470 373 6526
rect 175 6328 231 6384
rect 317 6328 373 6384
rect 175 6186 231 6242
rect 317 6186 373 6242
rect 175 6044 231 6100
rect 317 6044 373 6100
rect 175 5902 231 5958
rect 317 5902 373 5958
rect 175 5760 231 5816
rect 317 5760 373 5816
rect 175 5618 231 5674
rect 317 5618 373 5674
rect 175 5476 231 5532
rect 317 5476 373 5532
rect 175 5334 231 5390
rect 317 5334 373 5390
rect 175 5192 231 5248
rect 317 5192 373 5248
rect 175 5050 231 5106
rect 317 5050 373 5106
rect 175 4908 231 4964
rect 317 4908 373 4964
rect 175 4766 231 4822
rect 317 4766 373 4822
rect 175 4624 231 4680
rect 317 4624 373 4680
rect 175 4482 231 4538
rect 317 4482 373 4538
rect 175 4122 231 4178
rect 317 4122 373 4178
rect 175 3980 231 4036
rect 317 3980 373 4036
rect 175 3838 231 3894
rect 317 3838 373 3894
rect 175 3696 231 3752
rect 317 3696 373 3752
rect 175 3554 231 3610
rect 317 3554 373 3610
rect 175 3412 231 3468
rect 317 3412 373 3468
rect 175 3270 231 3326
rect 317 3270 373 3326
rect 175 3128 231 3184
rect 317 3128 373 3184
rect 175 2986 231 3042
rect 317 2986 373 3042
rect 175 2844 231 2900
rect 317 2844 373 2900
rect 175 2702 231 2758
rect 317 2702 373 2758
rect 175 2560 231 2616
rect 317 2560 373 2616
rect 175 2418 231 2474
rect 317 2418 373 2474
rect 175 2276 231 2332
rect 317 2276 373 2332
rect 175 2134 231 2190
rect 317 2134 373 2190
rect 175 1992 231 2048
rect 317 1992 373 2048
rect 175 1850 231 1906
rect 317 1850 373 1906
rect 175 1708 231 1764
rect 317 1708 373 1764
rect 175 1566 231 1622
rect 317 1566 373 1622
rect 175 1424 231 1480
rect 317 1424 373 1480
rect 175 1282 231 1338
rect 317 1282 373 1338
<< metal3 >>
rect 1886 56865 1962 56875
rect 1886 56809 1896 56865
rect 1952 56809 1962 56865
rect 1886 56723 1962 56809
rect 1886 56667 1896 56723
rect 1952 56667 1962 56723
rect 1886 56581 1962 56667
rect 1886 56525 1896 56581
rect 1952 56525 1962 56581
rect 1886 56439 1962 56525
rect 2490 56810 13642 56820
rect 2490 56754 2500 56810
rect 2556 56754 2642 56810
rect 2698 56754 2784 56810
rect 2840 56754 2926 56810
rect 2982 56754 3068 56810
rect 3124 56754 3210 56810
rect 3266 56754 3352 56810
rect 3408 56754 3494 56810
rect 3550 56754 3636 56810
rect 3692 56754 3778 56810
rect 3834 56754 3920 56810
rect 3976 56754 4062 56810
rect 4118 56754 4204 56810
rect 4260 56754 4346 56810
rect 4402 56754 4488 56810
rect 4544 56754 4630 56810
rect 4686 56754 4772 56810
rect 4828 56754 4914 56810
rect 4970 56754 5056 56810
rect 5112 56754 5198 56810
rect 5254 56754 5340 56810
rect 5396 56754 5482 56810
rect 5538 56754 5624 56810
rect 5680 56754 5766 56810
rect 5822 56754 5908 56810
rect 5964 56754 6050 56810
rect 6106 56754 6192 56810
rect 6248 56754 6334 56810
rect 6390 56754 6476 56810
rect 6532 56754 6618 56810
rect 6674 56754 6760 56810
rect 6816 56754 6902 56810
rect 6958 56754 7044 56810
rect 7100 56754 7186 56810
rect 7242 56754 7328 56810
rect 7384 56754 7470 56810
rect 7526 56754 7612 56810
rect 7668 56754 7754 56810
rect 7810 56754 7896 56810
rect 7952 56754 8038 56810
rect 8094 56754 8180 56810
rect 8236 56754 8322 56810
rect 8378 56754 8464 56810
rect 8520 56754 8606 56810
rect 8662 56754 8748 56810
rect 8804 56754 8890 56810
rect 8946 56754 9032 56810
rect 9088 56754 9174 56810
rect 9230 56754 9316 56810
rect 9372 56754 9458 56810
rect 9514 56754 9600 56810
rect 9656 56754 9742 56810
rect 9798 56754 9884 56810
rect 9940 56754 10026 56810
rect 10082 56754 10168 56810
rect 10224 56754 10310 56810
rect 10366 56754 10452 56810
rect 10508 56754 10594 56810
rect 10650 56754 10736 56810
rect 10792 56754 10878 56810
rect 10934 56754 11020 56810
rect 11076 56754 11162 56810
rect 11218 56754 11304 56810
rect 11360 56754 11446 56810
rect 11502 56754 11588 56810
rect 11644 56754 11730 56810
rect 11786 56754 11872 56810
rect 11928 56754 12014 56810
rect 12070 56754 12156 56810
rect 12212 56754 12298 56810
rect 12354 56754 12440 56810
rect 12496 56754 12582 56810
rect 12638 56754 12724 56810
rect 12780 56754 12866 56810
rect 12922 56754 13008 56810
rect 13064 56754 13150 56810
rect 13206 56754 13292 56810
rect 13348 56754 13434 56810
rect 13490 56754 13576 56810
rect 13632 56754 13642 56810
rect 2490 56668 13642 56754
rect 2490 56612 2500 56668
rect 2556 56612 2642 56668
rect 2698 56612 2784 56668
rect 2840 56612 2926 56668
rect 2982 56612 3068 56668
rect 3124 56612 3210 56668
rect 3266 56612 3352 56668
rect 3408 56612 3494 56668
rect 3550 56612 3636 56668
rect 3692 56612 3778 56668
rect 3834 56612 3920 56668
rect 3976 56612 4062 56668
rect 4118 56612 4204 56668
rect 4260 56612 4346 56668
rect 4402 56612 4488 56668
rect 4544 56612 4630 56668
rect 4686 56612 4772 56668
rect 4828 56612 4914 56668
rect 4970 56612 5056 56668
rect 5112 56612 5198 56668
rect 5254 56612 5340 56668
rect 5396 56612 5482 56668
rect 5538 56612 5624 56668
rect 5680 56612 5766 56668
rect 5822 56612 5908 56668
rect 5964 56612 6050 56668
rect 6106 56612 6192 56668
rect 6248 56612 6334 56668
rect 6390 56612 6476 56668
rect 6532 56612 6618 56668
rect 6674 56612 6760 56668
rect 6816 56612 6902 56668
rect 6958 56612 7044 56668
rect 7100 56612 7186 56668
rect 7242 56612 7328 56668
rect 7384 56612 7470 56668
rect 7526 56612 7612 56668
rect 7668 56612 7754 56668
rect 7810 56612 7896 56668
rect 7952 56612 8038 56668
rect 8094 56612 8180 56668
rect 8236 56612 8322 56668
rect 8378 56612 8464 56668
rect 8520 56612 8606 56668
rect 8662 56612 8748 56668
rect 8804 56612 8890 56668
rect 8946 56612 9032 56668
rect 9088 56612 9174 56668
rect 9230 56612 9316 56668
rect 9372 56612 9458 56668
rect 9514 56612 9600 56668
rect 9656 56612 9742 56668
rect 9798 56612 9884 56668
rect 9940 56612 10026 56668
rect 10082 56612 10168 56668
rect 10224 56612 10310 56668
rect 10366 56612 10452 56668
rect 10508 56612 10594 56668
rect 10650 56612 10736 56668
rect 10792 56612 10878 56668
rect 10934 56612 11020 56668
rect 11076 56612 11162 56668
rect 11218 56612 11304 56668
rect 11360 56612 11446 56668
rect 11502 56612 11588 56668
rect 11644 56612 11730 56668
rect 11786 56612 11872 56668
rect 11928 56612 12014 56668
rect 12070 56612 12156 56668
rect 12212 56612 12298 56668
rect 12354 56612 12440 56668
rect 12496 56612 12582 56668
rect 12638 56612 12724 56668
rect 12780 56612 12866 56668
rect 12922 56612 13008 56668
rect 13064 56612 13150 56668
rect 13206 56612 13292 56668
rect 13348 56612 13434 56668
rect 13490 56612 13576 56668
rect 13632 56612 13642 56668
rect 2490 56526 13642 56612
rect 2490 56470 2500 56526
rect 2556 56470 2642 56526
rect 2698 56470 2784 56526
rect 2840 56470 2926 56526
rect 2982 56470 3068 56526
rect 3124 56470 3210 56526
rect 3266 56470 3352 56526
rect 3408 56470 3494 56526
rect 3550 56470 3636 56526
rect 3692 56470 3778 56526
rect 3834 56470 3920 56526
rect 3976 56470 4062 56526
rect 4118 56470 4204 56526
rect 4260 56470 4346 56526
rect 4402 56470 4488 56526
rect 4544 56470 4630 56526
rect 4686 56470 4772 56526
rect 4828 56470 4914 56526
rect 4970 56470 5056 56526
rect 5112 56470 5198 56526
rect 5254 56470 5340 56526
rect 5396 56470 5482 56526
rect 5538 56470 5624 56526
rect 5680 56470 5766 56526
rect 5822 56470 5908 56526
rect 5964 56470 6050 56526
rect 6106 56470 6192 56526
rect 6248 56470 6334 56526
rect 6390 56470 6476 56526
rect 6532 56470 6618 56526
rect 6674 56470 6760 56526
rect 6816 56470 6902 56526
rect 6958 56470 7044 56526
rect 7100 56470 7186 56526
rect 7242 56470 7328 56526
rect 7384 56470 7470 56526
rect 7526 56470 7612 56526
rect 7668 56470 7754 56526
rect 7810 56470 7896 56526
rect 7952 56470 8038 56526
rect 8094 56470 8180 56526
rect 8236 56470 8322 56526
rect 8378 56470 8464 56526
rect 8520 56470 8606 56526
rect 8662 56470 8748 56526
rect 8804 56470 8890 56526
rect 8946 56470 9032 56526
rect 9088 56470 9174 56526
rect 9230 56470 9316 56526
rect 9372 56470 9458 56526
rect 9514 56470 9600 56526
rect 9656 56470 9742 56526
rect 9798 56470 9884 56526
rect 9940 56470 10026 56526
rect 10082 56470 10168 56526
rect 10224 56470 10310 56526
rect 10366 56470 10452 56526
rect 10508 56470 10594 56526
rect 10650 56470 10736 56526
rect 10792 56470 10878 56526
rect 10934 56470 11020 56526
rect 11076 56470 11162 56526
rect 11218 56470 11304 56526
rect 11360 56470 11446 56526
rect 11502 56470 11588 56526
rect 11644 56470 11730 56526
rect 11786 56470 11872 56526
rect 11928 56470 12014 56526
rect 12070 56470 12156 56526
rect 12212 56470 12298 56526
rect 12354 56470 12440 56526
rect 12496 56470 12582 56526
rect 12638 56470 12724 56526
rect 12780 56470 12866 56526
rect 12922 56470 13008 56526
rect 13064 56470 13150 56526
rect 13206 56470 13292 56526
rect 13348 56470 13434 56526
rect 13490 56470 13576 56526
rect 13632 56470 13642 56526
rect 2490 56460 13642 56470
rect 1886 56383 1896 56439
rect 1952 56383 1962 56439
rect 1886 56297 1962 56383
rect 1886 56241 1896 56297
rect 1952 56241 1962 56297
rect 1886 56155 1962 56241
rect 1886 56099 1896 56155
rect 1952 56099 1962 56155
rect 1886 56013 1962 56099
rect 1886 55957 1896 56013
rect 1952 55957 1962 56013
rect 1886 55871 1962 55957
rect 1886 55815 1896 55871
rect 1952 55815 1962 55871
rect 1886 55729 1962 55815
rect 1886 55673 1896 55729
rect 1952 55673 1962 55729
rect 2490 56068 13642 56078
rect 2490 56012 2500 56068
rect 2556 56012 2642 56068
rect 2698 56012 2784 56068
rect 2840 56012 2926 56068
rect 2982 56012 3068 56068
rect 3124 56012 3210 56068
rect 3266 56012 3352 56068
rect 3408 56012 3494 56068
rect 3550 56012 3636 56068
rect 3692 56012 3778 56068
rect 3834 56012 3920 56068
rect 3976 56012 4062 56068
rect 4118 56012 4204 56068
rect 4260 56012 4346 56068
rect 4402 56012 4488 56068
rect 4544 56012 4630 56068
rect 4686 56012 4772 56068
rect 4828 56012 4914 56068
rect 4970 56012 5056 56068
rect 5112 56012 5198 56068
rect 5254 56012 5340 56068
rect 5396 56012 5482 56068
rect 5538 56012 5624 56068
rect 5680 56012 5766 56068
rect 5822 56012 5908 56068
rect 5964 56012 6050 56068
rect 6106 56012 6192 56068
rect 6248 56012 6334 56068
rect 6390 56012 6476 56068
rect 6532 56012 6618 56068
rect 6674 56012 6760 56068
rect 6816 56012 6902 56068
rect 6958 56012 7044 56068
rect 7100 56012 7186 56068
rect 7242 56012 7328 56068
rect 7384 56012 7470 56068
rect 7526 56012 7612 56068
rect 7668 56012 7754 56068
rect 7810 56012 7896 56068
rect 7952 56012 8038 56068
rect 8094 56012 8180 56068
rect 8236 56012 8322 56068
rect 8378 56012 8464 56068
rect 8520 56012 8606 56068
rect 8662 56012 8748 56068
rect 8804 56012 8890 56068
rect 8946 56012 9032 56068
rect 9088 56012 9174 56068
rect 9230 56012 9316 56068
rect 9372 56012 9458 56068
rect 9514 56012 9600 56068
rect 9656 56012 9742 56068
rect 9798 56012 9884 56068
rect 9940 56012 10026 56068
rect 10082 56012 10168 56068
rect 10224 56012 10310 56068
rect 10366 56012 10452 56068
rect 10508 56012 10594 56068
rect 10650 56012 10736 56068
rect 10792 56012 10878 56068
rect 10934 56012 11020 56068
rect 11076 56012 11162 56068
rect 11218 56012 11304 56068
rect 11360 56012 11446 56068
rect 11502 56012 11588 56068
rect 11644 56012 11730 56068
rect 11786 56012 11872 56068
rect 11928 56012 12014 56068
rect 12070 56012 12156 56068
rect 12212 56012 12298 56068
rect 12354 56012 12440 56068
rect 12496 56012 12582 56068
rect 12638 56012 12724 56068
rect 12780 56012 12866 56068
rect 12922 56012 13008 56068
rect 13064 56012 13150 56068
rect 13206 56012 13292 56068
rect 13348 56012 13434 56068
rect 13490 56012 13576 56068
rect 13632 56012 13642 56068
rect 2490 55926 13642 56012
rect 2490 55870 2500 55926
rect 2556 55870 2642 55926
rect 2698 55870 2784 55926
rect 2840 55870 2926 55926
rect 2982 55870 3068 55926
rect 3124 55870 3210 55926
rect 3266 55870 3352 55926
rect 3408 55870 3494 55926
rect 3550 55870 3636 55926
rect 3692 55870 3778 55926
rect 3834 55870 3920 55926
rect 3976 55870 4062 55926
rect 4118 55870 4204 55926
rect 4260 55870 4346 55926
rect 4402 55870 4488 55926
rect 4544 55870 4630 55926
rect 4686 55870 4772 55926
rect 4828 55870 4914 55926
rect 4970 55870 5056 55926
rect 5112 55870 5198 55926
rect 5254 55870 5340 55926
rect 5396 55870 5482 55926
rect 5538 55870 5624 55926
rect 5680 55870 5766 55926
rect 5822 55870 5908 55926
rect 5964 55870 6050 55926
rect 6106 55870 6192 55926
rect 6248 55870 6334 55926
rect 6390 55870 6476 55926
rect 6532 55870 6618 55926
rect 6674 55870 6760 55926
rect 6816 55870 6902 55926
rect 6958 55870 7044 55926
rect 7100 55870 7186 55926
rect 7242 55870 7328 55926
rect 7384 55870 7470 55926
rect 7526 55870 7612 55926
rect 7668 55870 7754 55926
rect 7810 55870 7896 55926
rect 7952 55870 8038 55926
rect 8094 55870 8180 55926
rect 8236 55870 8322 55926
rect 8378 55870 8464 55926
rect 8520 55870 8606 55926
rect 8662 55870 8748 55926
rect 8804 55870 8890 55926
rect 8946 55870 9032 55926
rect 9088 55870 9174 55926
rect 9230 55870 9316 55926
rect 9372 55870 9458 55926
rect 9514 55870 9600 55926
rect 9656 55870 9742 55926
rect 9798 55870 9884 55926
rect 9940 55870 10026 55926
rect 10082 55870 10168 55926
rect 10224 55870 10310 55926
rect 10366 55870 10452 55926
rect 10508 55870 10594 55926
rect 10650 55870 10736 55926
rect 10792 55870 10878 55926
rect 10934 55870 11020 55926
rect 11076 55870 11162 55926
rect 11218 55870 11304 55926
rect 11360 55870 11446 55926
rect 11502 55870 11588 55926
rect 11644 55870 11730 55926
rect 11786 55870 11872 55926
rect 11928 55870 12014 55926
rect 12070 55870 12156 55926
rect 12212 55870 12298 55926
rect 12354 55870 12440 55926
rect 12496 55870 12582 55926
rect 12638 55870 12724 55926
rect 12780 55870 12866 55926
rect 12922 55870 13008 55926
rect 13064 55870 13150 55926
rect 13206 55870 13292 55926
rect 13348 55870 13434 55926
rect 13490 55870 13576 55926
rect 13632 55870 13642 55926
rect 2490 55784 13642 55870
rect 2490 55728 2500 55784
rect 2556 55728 2642 55784
rect 2698 55728 2784 55784
rect 2840 55728 2926 55784
rect 2982 55728 3068 55784
rect 3124 55728 3210 55784
rect 3266 55728 3352 55784
rect 3408 55728 3494 55784
rect 3550 55728 3636 55784
rect 3692 55728 3778 55784
rect 3834 55728 3920 55784
rect 3976 55728 4062 55784
rect 4118 55728 4204 55784
rect 4260 55728 4346 55784
rect 4402 55728 4488 55784
rect 4544 55728 4630 55784
rect 4686 55728 4772 55784
rect 4828 55728 4914 55784
rect 4970 55728 5056 55784
rect 5112 55728 5198 55784
rect 5254 55728 5340 55784
rect 5396 55728 5482 55784
rect 5538 55728 5624 55784
rect 5680 55728 5766 55784
rect 5822 55728 5908 55784
rect 5964 55728 6050 55784
rect 6106 55728 6192 55784
rect 6248 55728 6334 55784
rect 6390 55728 6476 55784
rect 6532 55728 6618 55784
rect 6674 55728 6760 55784
rect 6816 55728 6902 55784
rect 6958 55728 7044 55784
rect 7100 55728 7186 55784
rect 7242 55728 7328 55784
rect 7384 55728 7470 55784
rect 7526 55728 7612 55784
rect 7668 55728 7754 55784
rect 7810 55728 7896 55784
rect 7952 55728 8038 55784
rect 8094 55728 8180 55784
rect 8236 55728 8322 55784
rect 8378 55728 8464 55784
rect 8520 55728 8606 55784
rect 8662 55728 8748 55784
rect 8804 55728 8890 55784
rect 8946 55728 9032 55784
rect 9088 55728 9174 55784
rect 9230 55728 9316 55784
rect 9372 55728 9458 55784
rect 9514 55728 9600 55784
rect 9656 55728 9742 55784
rect 9798 55728 9884 55784
rect 9940 55728 10026 55784
rect 10082 55728 10168 55784
rect 10224 55728 10310 55784
rect 10366 55728 10452 55784
rect 10508 55728 10594 55784
rect 10650 55728 10736 55784
rect 10792 55728 10878 55784
rect 10934 55728 11020 55784
rect 11076 55728 11162 55784
rect 11218 55728 11304 55784
rect 11360 55728 11446 55784
rect 11502 55728 11588 55784
rect 11644 55728 11730 55784
rect 11786 55728 11872 55784
rect 11928 55728 12014 55784
rect 12070 55728 12156 55784
rect 12212 55728 12298 55784
rect 12354 55728 12440 55784
rect 12496 55728 12582 55784
rect 12638 55728 12724 55784
rect 12780 55728 12866 55784
rect 12922 55728 13008 55784
rect 13064 55728 13150 55784
rect 13206 55728 13292 55784
rect 13348 55728 13434 55784
rect 13490 55728 13576 55784
rect 13632 55728 13642 55784
rect 2490 55718 13642 55728
rect 1886 55663 1962 55673
rect 4758 55397 4834 55407
rect 4758 55341 4768 55397
rect 4824 55341 4834 55397
rect 4758 55255 4834 55341
rect 4758 55199 4768 55255
rect 4824 55199 4834 55255
rect 4758 55113 4834 55199
rect 4758 55057 4768 55113
rect 4824 55057 4834 55113
rect 4758 54971 4834 55057
rect 4758 54915 4768 54971
rect 4824 54915 4834 54971
rect 4758 54829 4834 54915
rect 4758 54773 4768 54829
rect 4824 54773 4834 54829
rect 4758 54687 4834 54773
rect 4758 54631 4768 54687
rect 4824 54631 4834 54687
rect 4758 54621 4834 54631
rect 4938 55397 5014 55407
rect 4938 55341 4948 55397
rect 5004 55341 5014 55397
rect 4938 55255 5014 55341
rect 4938 55199 4948 55255
rect 5004 55199 5014 55255
rect 4938 55113 5014 55199
rect 4938 55057 4948 55113
rect 5004 55057 5014 55113
rect 4938 54971 5014 55057
rect 4938 54915 4948 54971
rect 5004 54915 5014 54971
rect 4938 54829 5014 54915
rect 4938 54773 4948 54829
rect 5004 54773 5014 54829
rect 4938 54687 5014 54773
rect 4938 54631 4948 54687
rect 5004 54631 5014 54687
rect 4938 54621 5014 54631
rect 5426 55397 5502 55407
rect 5426 55341 5436 55397
rect 5492 55341 5502 55397
rect 5426 55255 5502 55341
rect 5426 55199 5436 55255
rect 5492 55199 5502 55255
rect 5426 55113 5502 55199
rect 5426 55057 5436 55113
rect 5492 55057 5502 55113
rect 5426 54971 5502 55057
rect 5426 54915 5436 54971
rect 5492 54915 5502 54971
rect 5426 54829 5502 54915
rect 5426 54773 5436 54829
rect 5492 54773 5502 54829
rect 5426 54687 5502 54773
rect 5426 54631 5436 54687
rect 5492 54631 5502 54687
rect 5426 54621 5502 54631
rect 5914 55397 5990 55407
rect 5914 55341 5924 55397
rect 5980 55341 5990 55397
rect 6278 55397 6354 55407
rect 5914 55255 5990 55341
rect 5914 55199 5924 55255
rect 5980 55199 5990 55255
rect 5914 55113 5990 55199
rect 5914 55057 5924 55113
rect 5980 55057 5990 55113
rect 5914 54971 5990 55057
rect 5914 54915 5924 54971
rect 5980 54915 5990 54971
rect 5914 54829 5990 54915
rect 5914 54773 5924 54829
rect 5980 54773 5990 54829
rect 5914 54687 5990 54773
rect 5914 54631 5924 54687
rect 5980 54631 5990 54687
rect 5914 54621 5990 54631
rect 6096 55371 6172 55381
rect 6096 55315 6106 55371
rect 6162 55315 6172 55371
rect 6096 55229 6172 55315
rect 6096 55173 6106 55229
rect 6162 55173 6172 55229
rect 6096 55087 6172 55173
rect 6096 55031 6106 55087
rect 6162 55031 6172 55087
rect 6096 54945 6172 55031
rect 6096 54889 6106 54945
rect 6162 54889 6172 54945
rect 6096 54803 6172 54889
rect 6096 54747 6106 54803
rect 6162 54747 6172 54803
rect 6096 54661 6172 54747
rect 6096 54605 6106 54661
rect 6162 54605 6172 54661
rect 6278 55341 6288 55397
rect 6344 55341 6354 55397
rect 6278 55255 6354 55341
rect 6278 55199 6288 55255
rect 6344 55199 6354 55255
rect 6278 55113 6354 55199
rect 6278 55057 6288 55113
rect 6344 55057 6354 55113
rect 6278 54971 6354 55057
rect 6278 54915 6288 54971
rect 6344 54915 6354 54971
rect 6278 54829 6354 54915
rect 6278 54773 6288 54829
rect 6344 54773 6354 54829
rect 6278 54687 6354 54773
rect 6278 54631 6288 54687
rect 6344 54631 6354 54687
rect 6278 54621 6354 54631
rect 6766 55397 6842 55407
rect 6766 55341 6776 55397
rect 6832 55341 6842 55397
rect 6766 55255 6842 55341
rect 6766 55199 6776 55255
rect 6832 55199 6842 55255
rect 6766 55113 6842 55199
rect 6766 55057 6776 55113
rect 6832 55057 6842 55113
rect 6766 54971 6842 55057
rect 6766 54915 6776 54971
rect 6832 54915 6842 54971
rect 6766 54829 6842 54915
rect 6766 54773 6776 54829
rect 6832 54773 6842 54829
rect 6766 54687 6842 54773
rect 6766 54631 6776 54687
rect 6832 54631 6842 54687
rect 6766 54621 6842 54631
rect 7254 55397 7330 55407
rect 7254 55341 7264 55397
rect 7320 55341 7330 55397
rect 7254 55255 7330 55341
rect 7254 55199 7264 55255
rect 7320 55199 7330 55255
rect 7254 55113 7330 55199
rect 7254 55057 7264 55113
rect 7320 55057 7330 55113
rect 7254 54971 7330 55057
rect 7254 54915 7264 54971
rect 7320 54915 7330 54971
rect 7254 54829 7330 54915
rect 7254 54773 7264 54829
rect 7320 54773 7330 54829
rect 7254 54687 7330 54773
rect 7254 54631 7264 54687
rect 7320 54631 7330 54687
rect 7254 54621 7330 54631
rect 7434 55397 7510 55407
rect 7434 55341 7444 55397
rect 7500 55341 7510 55397
rect 7434 55255 7510 55341
rect 7434 55199 7444 55255
rect 7500 55199 7510 55255
rect 7434 55113 7510 55199
rect 7434 55057 7444 55113
rect 7500 55057 7510 55113
rect 7434 54971 7510 55057
rect 7434 54915 7444 54971
rect 7500 54915 7510 54971
rect 7434 54829 7510 54915
rect 7434 54773 7444 54829
rect 7500 54773 7510 54829
rect 7434 54687 7510 54773
rect 7434 54631 7444 54687
rect 7500 54631 7510 54687
rect 7434 54621 7510 54631
rect 10002 55397 10078 55407
rect 10002 55341 10012 55397
rect 10068 55341 10078 55397
rect 10002 55255 10078 55341
rect 10002 55199 10012 55255
rect 10068 55199 10078 55255
rect 10002 55113 10078 55199
rect 10002 55057 10012 55113
rect 10068 55057 10078 55113
rect 10002 54971 10078 55057
rect 10002 54915 10012 54971
rect 10068 54915 10078 54971
rect 10002 54829 10078 54915
rect 10002 54773 10012 54829
rect 10068 54773 10078 54829
rect 10002 54687 10078 54773
rect 10002 54631 10012 54687
rect 10068 54631 10078 54687
rect 10002 54621 10078 54631
rect 10182 55397 10258 55407
rect 10182 55341 10192 55397
rect 10248 55341 10258 55397
rect 10182 55255 10258 55341
rect 10182 55199 10192 55255
rect 10248 55199 10258 55255
rect 10182 55113 10258 55199
rect 10182 55057 10192 55113
rect 10248 55057 10258 55113
rect 10182 54971 10258 55057
rect 10182 54915 10192 54971
rect 10248 54915 10258 54971
rect 10182 54829 10258 54915
rect 10182 54773 10192 54829
rect 10248 54773 10258 54829
rect 10182 54687 10258 54773
rect 10182 54631 10192 54687
rect 10248 54631 10258 54687
rect 10182 54621 10258 54631
rect 10670 55397 10746 55407
rect 10670 55341 10680 55397
rect 10736 55341 10746 55397
rect 10670 55255 10746 55341
rect 10670 55199 10680 55255
rect 10736 55199 10746 55255
rect 10670 55113 10746 55199
rect 10670 55057 10680 55113
rect 10736 55057 10746 55113
rect 10670 54971 10746 55057
rect 10670 54915 10680 54971
rect 10736 54915 10746 54971
rect 10670 54829 10746 54915
rect 10670 54773 10680 54829
rect 10736 54773 10746 54829
rect 10670 54687 10746 54773
rect 10670 54631 10680 54687
rect 10736 54631 10746 54687
rect 10670 54621 10746 54631
rect 11158 55397 11234 55407
rect 11158 55341 11168 55397
rect 11224 55341 11234 55397
rect 11522 55397 11598 55407
rect 11158 55255 11234 55341
rect 11158 55199 11168 55255
rect 11224 55199 11234 55255
rect 11158 55113 11234 55199
rect 11158 55057 11168 55113
rect 11224 55057 11234 55113
rect 11158 54971 11234 55057
rect 11158 54915 11168 54971
rect 11224 54915 11234 54971
rect 11158 54829 11234 54915
rect 11158 54773 11168 54829
rect 11224 54773 11234 54829
rect 11158 54687 11234 54773
rect 11158 54631 11168 54687
rect 11224 54631 11234 54687
rect 11158 54621 11234 54631
rect 11340 55371 11416 55381
rect 11340 55315 11350 55371
rect 11406 55315 11416 55371
rect 11340 55229 11416 55315
rect 11340 55173 11350 55229
rect 11406 55173 11416 55229
rect 11340 55087 11416 55173
rect 11340 55031 11350 55087
rect 11406 55031 11416 55087
rect 11340 54945 11416 55031
rect 11340 54889 11350 54945
rect 11406 54889 11416 54945
rect 11340 54803 11416 54889
rect 11340 54747 11350 54803
rect 11406 54747 11416 54803
rect 11340 54661 11416 54747
rect 6096 54519 6172 54605
rect 6096 54463 6106 54519
rect 6162 54463 6172 54519
rect 6096 54453 6172 54463
rect 11340 54605 11350 54661
rect 11406 54605 11416 54661
rect 11522 55341 11532 55397
rect 11588 55341 11598 55397
rect 11522 55255 11598 55341
rect 11522 55199 11532 55255
rect 11588 55199 11598 55255
rect 11522 55113 11598 55199
rect 11522 55057 11532 55113
rect 11588 55057 11598 55113
rect 11522 54971 11598 55057
rect 11522 54915 11532 54971
rect 11588 54915 11598 54971
rect 11522 54829 11598 54915
rect 11522 54773 11532 54829
rect 11588 54773 11598 54829
rect 11522 54687 11598 54773
rect 11522 54631 11532 54687
rect 11588 54631 11598 54687
rect 11522 54621 11598 54631
rect 12010 55397 12086 55407
rect 12010 55341 12020 55397
rect 12076 55341 12086 55397
rect 12010 55255 12086 55341
rect 12010 55199 12020 55255
rect 12076 55199 12086 55255
rect 12010 55113 12086 55199
rect 12010 55057 12020 55113
rect 12076 55057 12086 55113
rect 12010 54971 12086 55057
rect 12010 54915 12020 54971
rect 12076 54915 12086 54971
rect 12010 54829 12086 54915
rect 12010 54773 12020 54829
rect 12076 54773 12086 54829
rect 12010 54687 12086 54773
rect 12010 54631 12020 54687
rect 12076 54631 12086 54687
rect 12010 54621 12086 54631
rect 12498 55397 12574 55407
rect 12498 55341 12508 55397
rect 12564 55341 12574 55397
rect 12498 55255 12574 55341
rect 12498 55199 12508 55255
rect 12564 55199 12574 55255
rect 12498 55113 12574 55199
rect 12498 55057 12508 55113
rect 12564 55057 12574 55113
rect 12498 54971 12574 55057
rect 12498 54915 12508 54971
rect 12564 54915 12574 54971
rect 12498 54829 12574 54915
rect 12498 54773 12508 54829
rect 12564 54773 12574 54829
rect 12498 54687 12574 54773
rect 12498 54631 12508 54687
rect 12564 54631 12574 54687
rect 12498 54621 12574 54631
rect 12678 55397 12754 55407
rect 12678 55341 12688 55397
rect 12744 55341 12754 55397
rect 12678 55255 12754 55341
rect 12678 55199 12688 55255
rect 12744 55199 12754 55255
rect 12678 55113 12754 55199
rect 12678 55057 12688 55113
rect 12744 55057 12754 55113
rect 12678 54971 12754 55057
rect 12678 54915 12688 54971
rect 12744 54915 12754 54971
rect 12678 54829 12754 54915
rect 12678 54773 12688 54829
rect 12744 54773 12754 54829
rect 12678 54687 12754 54773
rect 12678 54631 12688 54687
rect 12744 54631 12754 54687
rect 12678 54621 12754 54631
rect 14400 55397 14760 55407
rect 14400 55341 14410 55397
rect 14466 55341 14552 55397
rect 14608 55341 14694 55397
rect 14750 55341 14760 55397
rect 14400 55255 14760 55341
rect 14400 55199 14410 55255
rect 14466 55199 14552 55255
rect 14608 55199 14694 55255
rect 14750 55199 14760 55255
rect 14400 55113 14760 55199
rect 14400 55057 14410 55113
rect 14466 55057 14552 55113
rect 14608 55057 14694 55113
rect 14750 55057 14760 55113
rect 14400 54971 14760 55057
rect 14400 54915 14410 54971
rect 14466 54915 14552 54971
rect 14608 54915 14694 54971
rect 14750 54915 14760 54971
rect 14400 54829 14760 54915
rect 14400 54773 14410 54829
rect 14466 54773 14552 54829
rect 14608 54773 14694 54829
rect 14750 54773 14760 54829
rect 14400 54687 14760 54773
rect 14400 54631 14410 54687
rect 14466 54631 14552 54687
rect 14608 54631 14694 54687
rect 14750 54631 14760 54687
rect 11340 54519 11416 54605
rect 11340 54463 11350 54519
rect 11406 54463 11416 54519
rect 11340 54453 11416 54463
rect 14400 54545 14760 54631
rect 14400 54489 14410 54545
rect 14466 54489 14552 54545
rect 14608 54489 14694 54545
rect 14750 54489 14760 54545
rect 14400 54403 14760 54489
rect 14400 54347 14410 54403
rect 14466 54347 14552 54403
rect 14608 54347 14694 54403
rect 14750 54347 14760 54403
rect 14400 54261 14760 54347
rect 14400 54205 14410 54261
rect 14466 54205 14552 54261
rect 14608 54205 14694 54261
rect 14750 54205 14760 54261
rect 14400 54119 14760 54205
rect 14400 54063 14410 54119
rect 14466 54063 14552 54119
rect 14608 54063 14694 54119
rect 14750 54063 14760 54119
rect 14400 54053 14760 54063
rect 6096 53814 6172 53824
rect 1886 53797 1962 53807
rect 1886 53741 1896 53797
rect 1952 53741 1962 53797
rect 1886 53655 1962 53741
rect 6096 53758 6106 53814
rect 6162 53758 6172 53814
rect 11340 53814 11416 53824
rect 1886 53599 1896 53655
rect 1952 53599 1962 53655
rect 1886 53513 1962 53599
rect 1886 53457 1896 53513
rect 1952 53457 1962 53513
rect 1886 53371 1962 53457
rect 1886 53315 1896 53371
rect 1952 53315 1962 53371
rect 1886 53229 1962 53315
rect 1886 53173 1896 53229
rect 1952 53173 1962 53229
rect 1886 53087 1962 53173
rect 1886 53031 1896 53087
rect 1952 53031 1962 53087
rect 1886 52945 1962 53031
rect 4758 53729 4834 53739
rect 4758 53673 4768 53729
rect 4824 53673 4834 53729
rect 4758 53587 4834 53673
rect 4758 53531 4768 53587
rect 4824 53531 4834 53587
rect 4758 53445 4834 53531
rect 4758 53389 4768 53445
rect 4824 53389 4834 53445
rect 4758 53303 4834 53389
rect 4758 53247 4768 53303
rect 4824 53247 4834 53303
rect 4758 53161 4834 53247
rect 4758 53105 4768 53161
rect 4824 53105 4834 53161
rect 4758 53019 4834 53105
rect 4758 52963 4768 53019
rect 4824 52963 4834 53019
rect 4758 52953 4834 52963
rect 4938 53729 5014 53739
rect 4938 53673 4948 53729
rect 5004 53673 5014 53729
rect 4938 53587 5014 53673
rect 4938 53531 4948 53587
rect 5004 53531 5014 53587
rect 4938 53445 5014 53531
rect 4938 53389 4948 53445
rect 5004 53389 5014 53445
rect 4938 53303 5014 53389
rect 4938 53247 4948 53303
rect 5004 53247 5014 53303
rect 4938 53161 5014 53247
rect 4938 53105 4948 53161
rect 5004 53105 5014 53161
rect 4938 53019 5014 53105
rect 4938 52963 4948 53019
rect 5004 52963 5014 53019
rect 4938 52953 5014 52963
rect 5426 53729 5502 53739
rect 5426 53673 5436 53729
rect 5492 53673 5502 53729
rect 5426 53587 5502 53673
rect 5426 53531 5436 53587
rect 5492 53531 5502 53587
rect 5426 53445 5502 53531
rect 5426 53389 5436 53445
rect 5492 53389 5502 53445
rect 5426 53303 5502 53389
rect 5426 53247 5436 53303
rect 5492 53247 5502 53303
rect 5426 53161 5502 53247
rect 5426 53105 5436 53161
rect 5492 53105 5502 53161
rect 5426 53019 5502 53105
rect 5426 52963 5436 53019
rect 5492 52963 5502 53019
rect 5426 52953 5502 52963
rect 5914 53729 5990 53739
rect 5914 53673 5924 53729
rect 5980 53673 5990 53729
rect 5914 53587 5990 53673
rect 5914 53531 5924 53587
rect 5980 53531 5990 53587
rect 5914 53445 5990 53531
rect 5914 53389 5924 53445
rect 5980 53389 5990 53445
rect 5914 53303 5990 53389
rect 5914 53247 5924 53303
rect 5980 53247 5990 53303
rect 5914 53161 5990 53247
rect 5914 53105 5924 53161
rect 5980 53105 5990 53161
rect 5914 53019 5990 53105
rect 5914 52963 5924 53019
rect 5980 52963 5990 53019
rect 5914 52953 5990 52963
rect 6096 53672 6172 53758
rect 9169 53797 9529 53807
rect 9169 53741 9179 53797
rect 9235 53741 9321 53797
rect 9377 53741 9463 53797
rect 9519 53741 9529 53797
rect 6096 53616 6106 53672
rect 6162 53616 6172 53672
rect 6096 53530 6172 53616
rect 6096 53474 6106 53530
rect 6162 53474 6172 53530
rect 6096 53388 6172 53474
rect 6096 53332 6106 53388
rect 6162 53332 6172 53388
rect 6096 53246 6172 53332
rect 6096 53190 6106 53246
rect 6162 53190 6172 53246
rect 6096 53104 6172 53190
rect 6096 53048 6106 53104
rect 6162 53048 6172 53104
rect 6096 52962 6172 53048
rect 1886 52889 1896 52945
rect 1952 52889 1962 52945
rect 6096 52906 6106 52962
rect 6162 52906 6172 52962
rect 6278 53729 6354 53739
rect 6278 53673 6288 53729
rect 6344 53673 6354 53729
rect 6278 53587 6354 53673
rect 6278 53531 6288 53587
rect 6344 53531 6354 53587
rect 6278 53445 6354 53531
rect 6278 53389 6288 53445
rect 6344 53389 6354 53445
rect 6278 53303 6354 53389
rect 6278 53247 6288 53303
rect 6344 53247 6354 53303
rect 6278 53161 6354 53247
rect 6278 53105 6288 53161
rect 6344 53105 6354 53161
rect 6278 53019 6354 53105
rect 6278 52963 6288 53019
rect 6344 52963 6354 53019
rect 6278 52953 6354 52963
rect 6766 53729 6842 53739
rect 6766 53673 6776 53729
rect 6832 53673 6842 53729
rect 6766 53587 6842 53673
rect 6766 53531 6776 53587
rect 6832 53531 6842 53587
rect 6766 53445 6842 53531
rect 6766 53389 6776 53445
rect 6832 53389 6842 53445
rect 6766 53303 6842 53389
rect 6766 53247 6776 53303
rect 6832 53247 6842 53303
rect 6766 53161 6842 53247
rect 6766 53105 6776 53161
rect 6832 53105 6842 53161
rect 6766 53019 6842 53105
rect 6766 52963 6776 53019
rect 6832 52963 6842 53019
rect 6766 52953 6842 52963
rect 7254 53729 7330 53739
rect 7254 53673 7264 53729
rect 7320 53673 7330 53729
rect 7254 53587 7330 53673
rect 7254 53531 7264 53587
rect 7320 53531 7330 53587
rect 7254 53445 7330 53531
rect 7254 53389 7264 53445
rect 7320 53389 7330 53445
rect 7254 53303 7330 53389
rect 7254 53247 7264 53303
rect 7320 53247 7330 53303
rect 7254 53161 7330 53247
rect 7254 53105 7264 53161
rect 7320 53105 7330 53161
rect 7254 53019 7330 53105
rect 7254 52963 7264 53019
rect 7320 52963 7330 53019
rect 7254 52953 7330 52963
rect 7434 53729 7510 53739
rect 7434 53673 7444 53729
rect 7500 53673 7510 53729
rect 7434 53587 7510 53673
rect 7434 53531 7444 53587
rect 7500 53531 7510 53587
rect 7434 53445 7510 53531
rect 7434 53389 7444 53445
rect 7500 53389 7510 53445
rect 7434 53303 7510 53389
rect 7434 53247 7444 53303
rect 7500 53247 7510 53303
rect 7434 53161 7510 53247
rect 7434 53105 7444 53161
rect 7500 53105 7510 53161
rect 7434 53019 7510 53105
rect 7434 52963 7444 53019
rect 7500 52963 7510 53019
rect 7434 52953 7510 52963
rect 9169 53655 9529 53741
rect 11340 53758 11350 53814
rect 11406 53758 11416 53814
rect 9169 53599 9179 53655
rect 9235 53599 9321 53655
rect 9377 53599 9463 53655
rect 9519 53599 9529 53655
rect 9169 53513 9529 53599
rect 9169 53457 9179 53513
rect 9235 53457 9321 53513
rect 9377 53457 9463 53513
rect 9519 53457 9529 53513
rect 9169 53371 9529 53457
rect 9169 53315 9179 53371
rect 9235 53315 9321 53371
rect 9377 53315 9463 53371
rect 9519 53315 9529 53371
rect 9169 53229 9529 53315
rect 9169 53173 9179 53229
rect 9235 53173 9321 53229
rect 9377 53173 9463 53229
rect 9519 53173 9529 53229
rect 9169 53087 9529 53173
rect 9169 53031 9179 53087
rect 9235 53031 9321 53087
rect 9377 53031 9463 53087
rect 9519 53031 9529 53087
rect 6096 52896 6172 52906
rect 9169 52945 9529 53031
rect 10002 53729 10078 53739
rect 10002 53673 10012 53729
rect 10068 53673 10078 53729
rect 10002 53587 10078 53673
rect 10002 53531 10012 53587
rect 10068 53531 10078 53587
rect 10002 53445 10078 53531
rect 10002 53389 10012 53445
rect 10068 53389 10078 53445
rect 10002 53303 10078 53389
rect 10002 53247 10012 53303
rect 10068 53247 10078 53303
rect 10002 53161 10078 53247
rect 10002 53105 10012 53161
rect 10068 53105 10078 53161
rect 10002 53019 10078 53105
rect 10002 52963 10012 53019
rect 10068 52963 10078 53019
rect 10002 52953 10078 52963
rect 10182 53729 10258 53739
rect 10182 53673 10192 53729
rect 10248 53673 10258 53729
rect 10182 53587 10258 53673
rect 10182 53531 10192 53587
rect 10248 53531 10258 53587
rect 10182 53445 10258 53531
rect 10182 53389 10192 53445
rect 10248 53389 10258 53445
rect 10182 53303 10258 53389
rect 10182 53247 10192 53303
rect 10248 53247 10258 53303
rect 10182 53161 10258 53247
rect 10182 53105 10192 53161
rect 10248 53105 10258 53161
rect 10182 53019 10258 53105
rect 10182 52963 10192 53019
rect 10248 52963 10258 53019
rect 10182 52953 10258 52963
rect 10670 53729 10746 53739
rect 10670 53673 10680 53729
rect 10736 53673 10746 53729
rect 10670 53587 10746 53673
rect 10670 53531 10680 53587
rect 10736 53531 10746 53587
rect 10670 53445 10746 53531
rect 10670 53389 10680 53445
rect 10736 53389 10746 53445
rect 10670 53303 10746 53389
rect 10670 53247 10680 53303
rect 10736 53247 10746 53303
rect 10670 53161 10746 53247
rect 10670 53105 10680 53161
rect 10736 53105 10746 53161
rect 10670 53019 10746 53105
rect 10670 52963 10680 53019
rect 10736 52963 10746 53019
rect 10670 52953 10746 52963
rect 11158 53729 11234 53739
rect 11158 53673 11168 53729
rect 11224 53673 11234 53729
rect 11158 53587 11234 53673
rect 11158 53531 11168 53587
rect 11224 53531 11234 53587
rect 11158 53445 11234 53531
rect 11158 53389 11168 53445
rect 11224 53389 11234 53445
rect 11158 53303 11234 53389
rect 11158 53247 11168 53303
rect 11224 53247 11234 53303
rect 11158 53161 11234 53247
rect 11158 53105 11168 53161
rect 11224 53105 11234 53161
rect 11158 53019 11234 53105
rect 11158 52963 11168 53019
rect 11224 52963 11234 53019
rect 11158 52953 11234 52963
rect 11340 53672 11416 53758
rect 11340 53616 11350 53672
rect 11406 53616 11416 53672
rect 11340 53530 11416 53616
rect 11340 53474 11350 53530
rect 11406 53474 11416 53530
rect 11340 53388 11416 53474
rect 11340 53332 11350 53388
rect 11406 53332 11416 53388
rect 11340 53246 11416 53332
rect 11340 53190 11350 53246
rect 11406 53190 11416 53246
rect 11340 53104 11416 53190
rect 11340 53048 11350 53104
rect 11406 53048 11416 53104
rect 11340 52962 11416 53048
rect 1886 52803 1962 52889
rect 1886 52747 1896 52803
rect 1952 52747 1962 52803
rect 1886 52661 1962 52747
rect 1886 52605 1896 52661
rect 1952 52605 1962 52661
rect 1886 52519 1962 52605
rect 1886 52463 1896 52519
rect 1952 52463 1962 52519
rect 1886 52453 1962 52463
rect 9169 52889 9179 52945
rect 9235 52889 9321 52945
rect 9377 52889 9463 52945
rect 9519 52889 9529 52945
rect 11340 52906 11350 52962
rect 11406 52906 11416 52962
rect 11522 53729 11598 53739
rect 11522 53673 11532 53729
rect 11588 53673 11598 53729
rect 11522 53587 11598 53673
rect 11522 53531 11532 53587
rect 11588 53531 11598 53587
rect 11522 53445 11598 53531
rect 11522 53389 11532 53445
rect 11588 53389 11598 53445
rect 11522 53303 11598 53389
rect 11522 53247 11532 53303
rect 11588 53247 11598 53303
rect 11522 53161 11598 53247
rect 11522 53105 11532 53161
rect 11588 53105 11598 53161
rect 11522 53019 11598 53105
rect 11522 52963 11532 53019
rect 11588 52963 11598 53019
rect 11522 52953 11598 52963
rect 12010 53729 12086 53739
rect 12010 53673 12020 53729
rect 12076 53673 12086 53729
rect 12010 53587 12086 53673
rect 12010 53531 12020 53587
rect 12076 53531 12086 53587
rect 12010 53445 12086 53531
rect 12010 53389 12020 53445
rect 12076 53389 12086 53445
rect 12010 53303 12086 53389
rect 12010 53247 12020 53303
rect 12076 53247 12086 53303
rect 12010 53161 12086 53247
rect 12010 53105 12020 53161
rect 12076 53105 12086 53161
rect 12010 53019 12086 53105
rect 12010 52963 12020 53019
rect 12076 52963 12086 53019
rect 12010 52953 12086 52963
rect 12498 53729 12574 53739
rect 12498 53673 12508 53729
rect 12564 53673 12574 53729
rect 12498 53587 12574 53673
rect 12498 53531 12508 53587
rect 12564 53531 12574 53587
rect 12498 53445 12574 53531
rect 12498 53389 12508 53445
rect 12564 53389 12574 53445
rect 12498 53303 12574 53389
rect 12498 53247 12508 53303
rect 12564 53247 12574 53303
rect 12498 53161 12574 53247
rect 12498 53105 12508 53161
rect 12564 53105 12574 53161
rect 12498 53019 12574 53105
rect 12498 52963 12508 53019
rect 12564 52963 12574 53019
rect 12498 52953 12574 52963
rect 12678 53729 12754 53739
rect 12678 53673 12688 53729
rect 12744 53673 12754 53729
rect 12678 53587 12754 53673
rect 12678 53531 12688 53587
rect 12744 53531 12754 53587
rect 12678 53445 12754 53531
rect 12678 53389 12688 53445
rect 12744 53389 12754 53445
rect 12678 53303 12754 53389
rect 12678 53247 12688 53303
rect 12744 53247 12754 53303
rect 12678 53161 12754 53247
rect 12678 53105 12688 53161
rect 12744 53105 12754 53161
rect 12678 53019 12754 53105
rect 12678 52963 12688 53019
rect 12744 52963 12754 53019
rect 12678 52953 12754 52963
rect 11340 52896 11416 52906
rect 9169 52803 9529 52889
rect 9169 52747 9179 52803
rect 9235 52747 9321 52803
rect 9377 52747 9463 52803
rect 9519 52747 9529 52803
rect 9169 52661 9529 52747
rect 9169 52605 9179 52661
rect 9235 52605 9321 52661
rect 9377 52605 9463 52661
rect 9519 52605 9529 52661
rect 9169 52519 9529 52605
rect 9169 52463 9179 52519
rect 9235 52463 9321 52519
rect 9377 52463 9463 52519
rect 9519 52463 9529 52519
rect 9169 52453 9529 52463
rect 46 52197 122 52207
rect 46 52141 56 52197
rect 112 52141 122 52197
rect 46 52055 122 52141
rect 46 51999 56 52055
rect 112 51999 122 52055
rect 46 51913 122 51999
rect 46 51857 56 51913
rect 112 51857 122 51913
rect 46 51771 122 51857
rect 46 51715 56 51771
rect 112 51715 122 51771
rect 46 51629 122 51715
rect 46 51573 56 51629
rect 112 51573 122 51629
rect 46 51487 122 51573
rect 46 51431 56 51487
rect 112 51431 122 51487
rect 46 51345 122 51431
rect 46 51289 56 51345
rect 112 51289 122 51345
rect 46 51203 122 51289
rect 46 51147 56 51203
rect 112 51147 122 51203
rect 46 51061 122 51147
rect 46 51005 56 51061
rect 112 51005 122 51061
rect 46 50919 122 51005
rect 46 50863 56 50919
rect 112 50863 122 50919
rect 46 50853 122 50863
rect 724 52197 1084 52207
rect 724 52141 734 52197
rect 790 52141 876 52197
rect 932 52141 1018 52197
rect 1074 52141 1084 52197
rect 724 52055 1084 52141
rect 724 51999 734 52055
rect 790 51999 876 52055
rect 932 51999 1018 52055
rect 1074 51999 1084 52055
rect 724 51913 1084 51999
rect 724 51857 734 51913
rect 790 51857 876 51913
rect 932 51857 1018 51913
rect 1074 51857 1084 51913
rect 724 51771 1084 51857
rect 724 51715 734 51771
rect 790 51715 876 51771
rect 932 51715 1018 51771
rect 1074 51715 1084 51771
rect 724 51629 1084 51715
rect 724 51573 734 51629
rect 790 51573 876 51629
rect 932 51573 1018 51629
rect 1074 51573 1084 51629
rect 724 51487 1084 51573
rect 724 51431 734 51487
rect 790 51431 876 51487
rect 932 51431 1018 51487
rect 1074 51431 1084 51487
rect 724 51345 1084 51431
rect 724 51289 734 51345
rect 790 51289 876 51345
rect 932 51289 1018 51345
rect 1074 51289 1084 51345
rect 724 51203 1084 51289
rect 724 51147 734 51203
rect 790 51147 876 51203
rect 932 51147 1018 51203
rect 1074 51147 1084 51203
rect 724 51061 1084 51147
rect 724 51005 734 51061
rect 790 51005 876 51061
rect 932 51005 1018 51061
rect 1074 51005 1084 51061
rect 724 50919 1084 51005
rect 724 50863 734 50919
rect 790 50863 876 50919
rect 932 50863 1018 50919
rect 1074 50863 1084 50919
rect 724 50853 1084 50863
rect 14942 52197 15018 52207
rect 14942 52141 14952 52197
rect 15008 52141 15018 52197
rect 14942 52055 15018 52141
rect 14942 51999 14952 52055
rect 15008 51999 15018 52055
rect 14942 51913 15018 51999
rect 14942 51857 14952 51913
rect 15008 51857 15018 51913
rect 14942 51771 15018 51857
rect 14942 51715 14952 51771
rect 15008 51715 15018 51771
rect 14942 51629 15018 51715
rect 14942 51573 14952 51629
rect 15008 51573 15018 51629
rect 14942 51487 15018 51573
rect 14942 51431 14952 51487
rect 15008 51431 15018 51487
rect 14942 51345 15018 51431
rect 14942 51289 14952 51345
rect 15008 51289 15018 51345
rect 14942 51203 15018 51289
rect 14942 51147 14952 51203
rect 15008 51147 15018 51203
rect 14942 51061 15018 51147
rect 14942 51005 14952 51061
rect 15008 51005 15018 51061
rect 14942 50919 15018 51005
rect 14942 50863 14952 50919
rect 15008 50863 15018 50919
rect 14942 50853 15018 50863
rect 204 50597 564 50607
rect 204 50541 214 50597
rect 270 50541 356 50597
rect 412 50541 498 50597
rect 554 50541 564 50597
rect 204 50455 564 50541
rect 204 50399 214 50455
rect 270 50399 356 50455
rect 412 50399 498 50455
rect 554 50399 564 50455
rect 204 50313 564 50399
rect 204 50257 214 50313
rect 270 50257 356 50313
rect 412 50257 498 50313
rect 554 50257 564 50313
rect 204 50171 564 50257
rect 204 50115 214 50171
rect 270 50115 356 50171
rect 412 50115 498 50171
rect 554 50115 564 50171
rect 204 50029 564 50115
rect 204 49973 214 50029
rect 270 49973 356 50029
rect 412 49973 498 50029
rect 554 49973 564 50029
rect 204 49887 564 49973
rect 204 49831 214 49887
rect 270 49831 356 49887
rect 412 49831 498 49887
rect 554 49831 564 49887
rect 204 49745 564 49831
rect 204 49689 214 49745
rect 270 49689 356 49745
rect 412 49689 498 49745
rect 554 49689 564 49745
rect 204 49603 564 49689
rect 204 49547 214 49603
rect 270 49547 356 49603
rect 412 49547 498 49603
rect 554 49547 564 49603
rect 204 49461 564 49547
rect 204 49405 214 49461
rect 270 49405 356 49461
rect 412 49405 498 49461
rect 554 49405 564 49461
rect 204 49319 564 49405
rect 204 49263 214 49319
rect 270 49263 356 49319
rect 412 49263 498 49319
rect 554 49263 564 49319
rect 11552 49568 11740 49578
rect 11552 49512 11562 49568
rect 11618 49512 11674 49568
rect 11730 49512 11740 49568
rect 11552 49456 11740 49512
rect 11552 49400 11562 49456
rect 11618 49400 11674 49456
rect 11730 49400 11740 49456
rect 11552 49344 11740 49400
rect 11552 49288 11562 49344
rect 11618 49288 11674 49344
rect 11730 49288 11740 49344
rect 11552 49278 11740 49288
rect 204 49253 564 49263
rect 10782 49014 10858 49024
rect 10782 48958 10792 49014
rect 10848 48958 10858 49014
rect 3978 48918 4302 48928
rect 3978 48862 3988 48918
rect 4044 48862 4112 48918
rect 4168 48862 4236 48918
rect 4292 48862 4302 48918
rect 3978 48794 4302 48862
rect 3978 48738 3988 48794
rect 4044 48738 4112 48794
rect 4168 48738 4236 48794
rect 4292 48738 4302 48794
rect 3978 48670 4302 48738
rect 3978 48614 3988 48670
rect 4044 48614 4112 48670
rect 4168 48614 4236 48670
rect 4292 48614 4302 48670
rect 3978 48546 4302 48614
rect 3978 48490 3988 48546
rect 4044 48490 4112 48546
rect 4168 48490 4236 48546
rect 4292 48490 4302 48546
rect 3978 48422 4302 48490
rect 3978 48366 3988 48422
rect 4044 48366 4112 48422
rect 4168 48366 4236 48422
rect 4292 48366 4302 48422
rect 3978 48298 4302 48366
rect 3978 48242 3988 48298
rect 4044 48242 4112 48298
rect 4168 48242 4236 48298
rect 4292 48242 4302 48298
rect 3978 48174 4302 48242
rect 3978 48118 3988 48174
rect 4044 48118 4112 48174
rect 4168 48118 4236 48174
rect 4292 48118 4302 48174
rect 3978 48050 4302 48118
rect 3978 47994 3988 48050
rect 4044 47994 4112 48050
rect 4168 47994 4236 48050
rect 4292 47994 4302 48050
rect 3978 47926 4302 47994
rect 10782 48872 10858 48958
rect 10782 48816 10792 48872
rect 10848 48816 10858 48872
rect 10782 48730 10858 48816
rect 10782 48674 10792 48730
rect 10848 48674 10858 48730
rect 10782 48588 10858 48674
rect 10782 48532 10792 48588
rect 10848 48532 10858 48588
rect 10782 48446 10858 48532
rect 10782 48390 10792 48446
rect 10848 48390 10858 48446
rect 10782 48304 10858 48390
rect 10782 48248 10792 48304
rect 10848 48248 10858 48304
rect 10782 48162 10858 48248
rect 10782 48106 10792 48162
rect 10848 48106 10858 48162
rect 10782 48020 10858 48106
rect 10782 47964 10792 48020
rect 10848 47964 10858 48020
rect 10782 47954 10858 47964
rect 3978 47870 3988 47926
rect 4044 47870 4112 47926
rect 4168 47870 4236 47926
rect 4292 47870 4302 47926
rect 3978 47802 4302 47870
rect 3978 47746 3988 47802
rect 4044 47746 4112 47802
rect 4168 47746 4236 47802
rect 4292 47746 4302 47802
rect 3978 47736 4302 47746
rect 3608 47414 3684 47424
rect 3608 47358 3618 47414
rect 3674 47358 3684 47414
rect 3608 47272 3684 47358
rect 3608 47216 3618 47272
rect 3674 47216 3684 47272
rect 3608 47130 3684 47216
rect 3608 47074 3618 47130
rect 3674 47074 3684 47130
rect 3608 46988 3684 47074
rect 3608 46932 3618 46988
rect 3674 46932 3684 46988
rect 3608 46846 3684 46932
rect 3608 46790 3618 46846
rect 3674 46790 3684 46846
rect 3608 46704 3684 46790
rect 3608 46648 3618 46704
rect 3674 46648 3684 46704
rect 3608 46562 3684 46648
rect 11001 47397 11077 47407
rect 11001 47341 11011 47397
rect 11067 47341 11077 47397
rect 11001 47255 11077 47341
rect 11001 47199 11011 47255
rect 11067 47199 11077 47255
rect 11001 47113 11077 47199
rect 11001 47057 11011 47113
rect 11067 47057 11077 47113
rect 11001 46971 11077 47057
rect 11001 46915 11011 46971
rect 11067 46915 11077 46971
rect 11001 46829 11077 46915
rect 11001 46773 11011 46829
rect 11067 46773 11077 46829
rect 11001 46687 11077 46773
rect 11001 46631 11011 46687
rect 11067 46631 11077 46687
rect 11001 46621 11077 46631
rect 3608 46506 3618 46562
rect 3674 46506 3684 46562
rect 3608 46420 3684 46506
rect 3608 46364 3618 46420
rect 3674 46364 3684 46420
rect 3608 46354 3684 46364
rect 3969 45341 4293 45351
rect 3969 45285 3979 45341
rect 4035 45285 4103 45341
rect 4159 45285 4227 45341
rect 4283 45285 4293 45341
rect 3969 45217 4293 45285
rect 3969 45161 3979 45217
rect 4035 45161 4103 45217
rect 4159 45161 4227 45217
rect 4283 45161 4293 45217
rect 3969 45093 4293 45161
rect 3969 45037 3979 45093
rect 4035 45037 4103 45093
rect 4159 45037 4227 45093
rect 4283 45037 4293 45093
rect 3969 44969 4293 45037
rect 3969 44913 3979 44969
rect 4035 44913 4103 44969
rect 4159 44913 4227 44969
rect 4283 44913 4293 44969
rect 3969 44845 4293 44913
rect 3969 44789 3979 44845
rect 4035 44789 4103 44845
rect 4159 44789 4227 44845
rect 4283 44789 4293 44845
rect 3969 44721 4293 44789
rect 3969 44665 3979 44721
rect 4035 44665 4103 44721
rect 4159 44665 4227 44721
rect 4283 44665 4293 44721
rect 3969 44597 4293 44665
rect 3969 44541 3979 44597
rect 4035 44541 4103 44597
rect 4159 44541 4227 44597
rect 4283 44541 4293 44597
rect 3969 44531 4293 44541
rect 3608 44197 3684 44207
rect 3608 44141 3618 44197
rect 3674 44141 3684 44197
rect 3608 44055 3684 44141
rect 3608 43999 3618 44055
rect 3674 43999 3684 44055
rect 3608 43913 3684 43999
rect 3608 43857 3618 43913
rect 3674 43857 3684 43913
rect 3608 43771 3684 43857
rect 3608 43715 3618 43771
rect 3674 43715 3684 43771
rect 3608 43629 3684 43715
rect 3608 43573 3618 43629
rect 3674 43573 3684 43629
rect 3608 43487 3684 43573
rect 3608 43431 3618 43487
rect 3674 43431 3684 43487
rect 3608 43345 3684 43431
rect 3608 43289 3618 43345
rect 3674 43289 3684 43345
rect 3608 43203 3684 43289
rect 3608 43147 3618 43203
rect 3674 43147 3684 43203
rect 3608 43061 3684 43147
rect 3608 43005 3618 43061
rect 3674 43005 3684 43061
rect 3608 42919 3684 43005
rect 3608 42863 3618 42919
rect 3674 42863 3684 42919
rect 3608 42853 3684 42863
rect 14400 44197 14760 44207
rect 14400 44141 14410 44197
rect 14466 44141 14552 44197
rect 14608 44141 14694 44197
rect 14750 44141 14760 44197
rect 14400 44055 14760 44141
rect 14400 43999 14410 44055
rect 14466 43999 14552 44055
rect 14608 43999 14694 44055
rect 14750 43999 14760 44055
rect 14400 43913 14760 43999
rect 14400 43857 14410 43913
rect 14466 43857 14552 43913
rect 14608 43857 14694 43913
rect 14750 43857 14760 43913
rect 14400 43771 14760 43857
rect 14400 43715 14410 43771
rect 14466 43715 14552 43771
rect 14608 43715 14694 43771
rect 14750 43715 14760 43771
rect 14400 43629 14760 43715
rect 14400 43573 14410 43629
rect 14466 43573 14552 43629
rect 14608 43573 14694 43629
rect 14750 43573 14760 43629
rect 14400 43487 14760 43573
rect 14400 43431 14410 43487
rect 14466 43431 14552 43487
rect 14608 43431 14694 43487
rect 14750 43431 14760 43487
rect 14400 43345 14760 43431
rect 14400 43289 14410 43345
rect 14466 43289 14552 43345
rect 14608 43289 14694 43345
rect 14750 43289 14760 43345
rect 14400 43203 14760 43289
rect 14400 43147 14410 43203
rect 14466 43147 14552 43203
rect 14608 43147 14694 43203
rect 14750 43147 14760 43203
rect 14400 43061 14760 43147
rect 14400 43005 14410 43061
rect 14466 43005 14552 43061
rect 14608 43005 14694 43061
rect 14750 43005 14760 43061
rect 14400 42919 14760 43005
rect 14400 42863 14410 42919
rect 14466 42863 14552 42919
rect 14608 42863 14694 42919
rect 14750 42863 14760 42919
rect 14400 42853 14760 42863
rect 3608 42597 3684 42607
rect 3608 42541 3618 42597
rect 3674 42541 3684 42597
rect 3608 42455 3684 42541
rect 3608 42399 3618 42455
rect 3674 42399 3684 42455
rect 3608 42313 3684 42399
rect 3608 42257 3618 42313
rect 3674 42257 3684 42313
rect 3608 42171 3684 42257
rect 3608 42115 3618 42171
rect 3674 42115 3684 42171
rect 3608 42029 3684 42115
rect 3608 41973 3618 42029
rect 3674 41973 3684 42029
rect 3608 41887 3684 41973
rect 3608 41831 3618 41887
rect 3674 41831 3684 41887
rect 3608 41745 3684 41831
rect 3608 41689 3618 41745
rect 3674 41689 3684 41745
rect 3608 41603 3684 41689
rect 3608 41547 3618 41603
rect 3674 41547 3684 41603
rect 3608 41461 3684 41547
rect 3608 41405 3618 41461
rect 3674 41405 3684 41461
rect 13181 42598 13481 42608
rect 13181 42542 13191 42598
rect 13247 42542 13303 42598
rect 13359 42542 13415 42598
rect 13471 42542 13481 42598
rect 13181 42486 13481 42542
rect 13181 42430 13191 42486
rect 13247 42430 13303 42486
rect 13359 42430 13415 42486
rect 13471 42430 13481 42486
rect 13181 42374 13481 42430
rect 13181 42318 13191 42374
rect 13247 42318 13303 42374
rect 13359 42318 13415 42374
rect 13471 42318 13481 42374
rect 13181 42262 13481 42318
rect 13181 42206 13191 42262
rect 13247 42206 13303 42262
rect 13359 42206 13415 42262
rect 13471 42206 13481 42262
rect 13181 42150 13481 42206
rect 13181 42094 13191 42150
rect 13247 42094 13303 42150
rect 13359 42094 13415 42150
rect 13471 42094 13481 42150
rect 13181 42038 13481 42094
rect 13181 41982 13191 42038
rect 13247 41982 13303 42038
rect 13359 41982 13415 42038
rect 13471 41982 13481 42038
rect 13181 41926 13481 41982
rect 13181 41870 13191 41926
rect 13247 41870 13303 41926
rect 13359 41870 13415 41926
rect 13471 41870 13481 41926
rect 13181 41814 13481 41870
rect 13181 41758 13191 41814
rect 13247 41758 13303 41814
rect 13359 41758 13415 41814
rect 13471 41758 13481 41814
rect 13181 41702 13481 41758
rect 13181 41646 13191 41702
rect 13247 41646 13303 41702
rect 13359 41646 13415 41702
rect 13471 41646 13481 41702
rect 13181 41590 13481 41646
rect 13181 41534 13191 41590
rect 13247 41534 13303 41590
rect 13359 41534 13415 41590
rect 13471 41534 13481 41590
rect 13181 41478 13481 41534
rect 13181 41422 13191 41478
rect 13247 41422 13303 41478
rect 13359 41422 13415 41478
rect 13471 41422 13481 41478
rect 13181 41412 13481 41422
rect 14400 42597 14760 42607
rect 14400 42541 14410 42597
rect 14466 42541 14552 42597
rect 14608 42541 14694 42597
rect 14750 42541 14760 42597
rect 14400 42455 14760 42541
rect 14400 42399 14410 42455
rect 14466 42399 14552 42455
rect 14608 42399 14694 42455
rect 14750 42399 14760 42455
rect 14400 42313 14760 42399
rect 14400 42257 14410 42313
rect 14466 42257 14552 42313
rect 14608 42257 14694 42313
rect 14750 42257 14760 42313
rect 14400 42171 14760 42257
rect 14400 42115 14410 42171
rect 14466 42115 14552 42171
rect 14608 42115 14694 42171
rect 14750 42115 14760 42171
rect 14400 42029 14760 42115
rect 14400 41973 14410 42029
rect 14466 41973 14552 42029
rect 14608 41973 14694 42029
rect 14750 41973 14760 42029
rect 14400 41887 14760 41973
rect 14400 41831 14410 41887
rect 14466 41831 14552 41887
rect 14608 41831 14694 41887
rect 14750 41831 14760 41887
rect 14400 41745 14760 41831
rect 14400 41689 14410 41745
rect 14466 41689 14552 41745
rect 14608 41689 14694 41745
rect 14750 41689 14760 41745
rect 14400 41603 14760 41689
rect 14400 41547 14410 41603
rect 14466 41547 14552 41603
rect 14608 41547 14694 41603
rect 14750 41547 14760 41603
rect 14400 41461 14760 41547
rect 3608 41319 3684 41405
rect 3608 41263 3618 41319
rect 3674 41263 3684 41319
rect 3608 41253 3684 41263
rect 14400 41405 14410 41461
rect 14466 41405 14552 41461
rect 14608 41405 14694 41461
rect 14750 41405 14760 41461
rect 14400 41319 14760 41405
rect 14400 41263 14410 41319
rect 14466 41263 14552 41319
rect 14608 41263 14694 41319
rect 14750 41263 14760 41319
rect 14400 41253 14760 41263
rect 14400 40997 14760 41007
rect 14400 40941 14410 40997
rect 14466 40941 14552 40997
rect 14608 40941 14694 40997
rect 14750 40941 14760 40997
rect 14400 40855 14760 40941
rect 14400 40799 14410 40855
rect 14466 40799 14552 40855
rect 14608 40799 14694 40855
rect 14750 40799 14760 40855
rect 14400 40713 14760 40799
rect 1836 40702 3758 40712
rect 1836 40646 1846 40702
rect 1902 40646 1988 40702
rect 2044 40646 2130 40702
rect 2186 40646 2272 40702
rect 2328 40646 2414 40702
rect 2470 40646 2556 40702
rect 2612 40646 2698 40702
rect 2754 40646 2840 40702
rect 2896 40646 2982 40702
rect 3038 40646 3124 40702
rect 3180 40646 3266 40702
rect 3322 40646 3408 40702
rect 3464 40646 3550 40702
rect 3606 40646 3692 40702
rect 3748 40646 3758 40702
rect 1836 40636 3758 40646
rect 14400 40657 14410 40713
rect 14466 40657 14552 40713
rect 14608 40657 14694 40713
rect 14750 40657 14760 40713
rect 14400 40571 14760 40657
rect 14400 40515 14410 40571
rect 14466 40515 14552 40571
rect 14608 40515 14694 40571
rect 14750 40515 14760 40571
rect 14400 40429 14760 40515
rect 14400 40373 14410 40429
rect 14466 40373 14552 40429
rect 14608 40373 14694 40429
rect 14750 40373 14760 40429
rect 14400 40287 14760 40373
rect 14400 40231 14410 40287
rect 14466 40231 14552 40287
rect 14608 40231 14694 40287
rect 14750 40231 14760 40287
rect 14400 40145 14760 40231
rect 14400 40089 14410 40145
rect 14466 40089 14552 40145
rect 14608 40089 14694 40145
rect 14750 40089 14760 40145
rect 14400 40003 14760 40089
rect 2428 39946 4492 39956
rect 2428 39890 2438 39946
rect 2494 39890 2580 39946
rect 2636 39890 2722 39946
rect 2778 39890 2864 39946
rect 2920 39890 3006 39946
rect 3062 39890 3148 39946
rect 3204 39890 3290 39946
rect 3346 39890 3432 39946
rect 3488 39890 3574 39946
rect 3630 39890 3716 39946
rect 3772 39890 3858 39946
rect 3914 39890 4000 39946
rect 4056 39890 4142 39946
rect 4198 39890 4284 39946
rect 4340 39890 4426 39946
rect 4482 39890 4492 39946
rect 2428 39880 4492 39890
rect 7987 39946 9767 39956
rect 7987 39890 7997 39946
rect 8053 39890 8139 39946
rect 8195 39890 8281 39946
rect 8337 39890 8423 39946
rect 8479 39890 8565 39946
rect 8621 39890 8707 39946
rect 8763 39890 8849 39946
rect 8905 39890 8991 39946
rect 9047 39890 9133 39946
rect 9189 39890 9275 39946
rect 9331 39890 9417 39946
rect 9473 39890 9559 39946
rect 9615 39890 9701 39946
rect 9757 39890 9767 39946
rect 7987 39880 9767 39890
rect 12748 39946 13818 39956
rect 12748 39890 12758 39946
rect 12814 39890 12900 39946
rect 12956 39890 13042 39946
rect 13098 39890 13184 39946
rect 13240 39890 13326 39946
rect 13382 39890 13468 39946
rect 13524 39890 13610 39946
rect 13666 39890 13752 39946
rect 13808 39890 13818 39946
rect 12748 39880 13818 39890
rect 14400 39947 14410 40003
rect 14466 39947 14552 40003
rect 14608 39947 14694 40003
rect 14750 39947 14760 40003
rect 14400 39861 14760 39947
rect 14400 39805 14410 39861
rect 14466 39805 14552 39861
rect 14608 39805 14694 39861
rect 14750 39805 14760 39861
rect 14400 39719 14760 39805
rect 14400 39663 14410 39719
rect 14466 39663 14552 39719
rect 14608 39663 14694 39719
rect 14750 39663 14760 39719
rect 14400 39653 14760 39663
rect 1771 39420 1847 39430
rect 204 39397 564 39407
rect 204 39341 214 39397
rect 270 39341 356 39397
rect 412 39341 498 39397
rect 554 39341 564 39397
rect 204 39255 564 39341
rect 204 39199 214 39255
rect 270 39199 356 39255
rect 412 39199 498 39255
rect 554 39199 564 39255
rect 204 39113 564 39199
rect 204 39057 214 39113
rect 270 39057 356 39113
rect 412 39057 498 39113
rect 554 39057 564 39113
rect 204 38971 564 39057
rect 204 38915 214 38971
rect 270 38915 356 38971
rect 412 38915 498 38971
rect 554 38915 564 38971
rect 204 38829 564 38915
rect 204 38773 214 38829
rect 270 38773 356 38829
rect 412 38773 498 38829
rect 554 38773 564 38829
rect 1771 39364 1781 39420
rect 1837 39364 1847 39420
rect 1771 39278 1847 39364
rect 1771 39222 1781 39278
rect 1837 39222 1847 39278
rect 1771 39136 1847 39222
rect 1771 39080 1781 39136
rect 1837 39080 1847 39136
rect 1771 38994 1847 39080
rect 1771 38938 1781 38994
rect 1837 38938 1847 38994
rect 1771 38852 1847 38938
rect 1771 38796 1781 38852
rect 1837 38796 1847 38852
rect 1771 38786 1847 38796
rect 5083 39420 5159 39430
rect 5083 39364 5093 39420
rect 5149 39364 5159 39420
rect 5083 39278 5159 39364
rect 5083 39222 5093 39278
rect 5149 39222 5159 39278
rect 5083 39136 5159 39222
rect 5083 39080 5093 39136
rect 5149 39080 5159 39136
rect 5083 38994 5159 39080
rect 5083 38938 5093 38994
rect 5149 38938 5159 38994
rect 5083 38852 5159 38938
rect 5083 38796 5093 38852
rect 5149 38796 5159 38852
rect 5083 38786 5159 38796
rect 6049 39414 6125 39424
rect 6049 39358 6059 39414
rect 6115 39358 6125 39414
rect 6049 39272 6125 39358
rect 6049 39216 6059 39272
rect 6115 39216 6125 39272
rect 6049 39130 6125 39216
rect 6049 39074 6059 39130
rect 6115 39074 6125 39130
rect 6049 38988 6125 39074
rect 6049 38932 6059 38988
rect 6115 38932 6125 38988
rect 6049 38846 6125 38932
rect 6049 38790 6059 38846
rect 6115 38790 6125 38846
rect 204 38687 564 38773
rect 204 38631 214 38687
rect 270 38631 356 38687
rect 412 38631 498 38687
rect 554 38631 564 38687
rect 204 38545 564 38631
rect 204 38489 214 38545
rect 270 38489 356 38545
rect 412 38489 498 38545
rect 554 38489 564 38545
rect 204 38403 564 38489
rect 204 38347 214 38403
rect 270 38347 356 38403
rect 412 38347 498 38403
rect 554 38347 564 38403
rect 6049 38704 6125 38790
rect 7015 39420 7091 39430
rect 7015 39364 7025 39420
rect 7081 39364 7091 39420
rect 7015 39278 7091 39364
rect 7015 39222 7025 39278
rect 7081 39222 7091 39278
rect 7015 39136 7091 39222
rect 7015 39080 7025 39136
rect 7081 39080 7091 39136
rect 7015 38994 7091 39080
rect 7015 38938 7025 38994
rect 7081 38938 7091 38994
rect 7015 38852 7091 38938
rect 7015 38796 7025 38852
rect 7081 38796 7091 38852
rect 7015 38786 7091 38796
rect 10327 39414 10403 39424
rect 10327 39358 10337 39414
rect 10393 39358 10403 39414
rect 10327 39272 10403 39358
rect 10327 39216 10337 39272
rect 10393 39216 10403 39272
rect 10327 39130 10403 39216
rect 10327 39074 10337 39130
rect 10393 39074 10403 39130
rect 10327 38988 10403 39074
rect 10327 38932 10337 38988
rect 10393 38932 10403 38988
rect 10327 38846 10403 38932
rect 10327 38790 10337 38846
rect 10393 38790 10403 38846
rect 6049 38648 6059 38704
rect 6115 38648 6125 38704
rect 6049 38562 6125 38648
rect 6049 38506 6059 38562
rect 6115 38506 6125 38562
rect 6049 38420 6125 38506
rect 6049 38364 6059 38420
rect 6115 38364 6125 38420
rect 6049 38354 6125 38364
rect 10327 38704 10403 38790
rect 10327 38648 10337 38704
rect 10393 38648 10403 38704
rect 10327 38562 10403 38648
rect 10327 38506 10337 38562
rect 10393 38506 10403 38562
rect 10327 38420 10403 38506
rect 10327 38364 10337 38420
rect 10393 38364 10403 38420
rect 10327 38354 10403 38364
rect 11200 39414 11276 39424
rect 11200 39358 11210 39414
rect 11266 39358 11276 39414
rect 11200 39272 11276 39358
rect 11200 39216 11210 39272
rect 11266 39216 11276 39272
rect 11200 39130 11276 39216
rect 11200 39074 11210 39130
rect 11266 39074 11276 39130
rect 11200 38988 11276 39074
rect 11200 38932 11210 38988
rect 11266 38932 11276 38988
rect 11200 38846 11276 38932
rect 11200 38790 11210 38846
rect 11266 38790 11276 38846
rect 11200 38704 11276 38790
rect 11200 38648 11210 38704
rect 11266 38648 11276 38704
rect 11200 38562 11276 38648
rect 11200 38506 11210 38562
rect 11266 38506 11276 38562
rect 11200 38420 11276 38506
rect 11200 38364 11210 38420
rect 11266 38364 11276 38420
rect 11200 38354 11276 38364
rect 204 38261 564 38347
rect 204 38205 214 38261
rect 270 38205 356 38261
rect 412 38205 498 38261
rect 554 38205 564 38261
rect 204 38119 564 38205
rect 204 38063 214 38119
rect 270 38063 356 38119
rect 412 38063 498 38119
rect 554 38063 564 38119
rect 204 38053 564 38063
rect 46 37797 122 37807
rect 46 37741 56 37797
rect 112 37741 122 37797
rect 46 37655 122 37741
rect 46 37599 56 37655
rect 112 37599 122 37655
rect 46 37513 122 37599
rect 46 37457 56 37513
rect 112 37457 122 37513
rect 46 37371 122 37457
rect 46 37315 56 37371
rect 112 37315 122 37371
rect 46 37229 122 37315
rect 46 37173 56 37229
rect 112 37173 122 37229
rect 46 37087 122 37173
rect 46 37031 56 37087
rect 112 37031 122 37087
rect 46 36945 122 37031
rect 46 36889 56 36945
rect 112 36889 122 36945
rect 46 36803 122 36889
rect 46 36747 56 36803
rect 112 36747 122 36803
rect 46 36661 122 36747
rect 46 36605 56 36661
rect 112 36605 122 36661
rect 46 36519 122 36605
rect 46 36463 56 36519
rect 112 36463 122 36519
rect 46 36453 122 36463
rect 724 37797 1084 37807
rect 724 37741 734 37797
rect 790 37741 876 37797
rect 932 37741 1018 37797
rect 1074 37741 1084 37797
rect 724 37655 1084 37741
rect 724 37599 734 37655
rect 790 37599 876 37655
rect 932 37599 1018 37655
rect 1074 37599 1084 37655
rect 724 37513 1084 37599
rect 724 37457 734 37513
rect 790 37457 876 37513
rect 932 37457 1018 37513
rect 1074 37457 1084 37513
rect 724 37371 1084 37457
rect 724 37315 734 37371
rect 790 37315 876 37371
rect 932 37315 1018 37371
rect 1074 37315 1084 37371
rect 724 37229 1084 37315
rect 724 37173 734 37229
rect 790 37173 876 37229
rect 932 37173 1018 37229
rect 1074 37173 1084 37229
rect 724 37087 1084 37173
rect 724 37031 734 37087
rect 790 37031 876 37087
rect 932 37031 1018 37087
rect 1074 37031 1084 37087
rect 724 36945 1084 37031
rect 724 36889 734 36945
rect 790 36889 876 36945
rect 932 36889 1018 36945
rect 1074 36889 1084 36945
rect 724 36803 1084 36889
rect 724 36747 734 36803
rect 790 36747 876 36803
rect 932 36747 1018 36803
rect 1074 36747 1084 36803
rect 724 36661 1084 36747
rect 724 36605 734 36661
rect 790 36605 876 36661
rect 932 36605 1018 36661
rect 1074 36605 1084 36661
rect 724 36519 1084 36605
rect 724 36463 734 36519
rect 790 36463 876 36519
rect 932 36463 1018 36519
rect 1074 36463 1084 36519
rect 724 36453 1084 36463
rect 6049 37797 6125 37807
rect 6049 37741 6059 37797
rect 6115 37741 6125 37797
rect 6049 37655 6125 37741
rect 6049 37599 6059 37655
rect 6115 37599 6125 37655
rect 6049 37513 6125 37599
rect 6049 37457 6059 37513
rect 6115 37457 6125 37513
rect 6049 37371 6125 37457
rect 6049 37315 6059 37371
rect 6115 37315 6125 37371
rect 6049 37229 6125 37315
rect 6049 37173 6059 37229
rect 6115 37173 6125 37229
rect 12406 37797 12624 37807
rect 12406 37741 12416 37797
rect 12472 37741 12558 37797
rect 12614 37741 12624 37797
rect 12406 37655 12624 37741
rect 12406 37599 12416 37655
rect 12472 37599 12558 37655
rect 12614 37599 12624 37655
rect 12406 37513 12624 37599
rect 12406 37457 12416 37513
rect 12472 37457 12558 37513
rect 12614 37457 12624 37513
rect 12406 37371 12624 37457
rect 12406 37315 12416 37371
rect 12472 37315 12558 37371
rect 12614 37315 12624 37371
rect 12406 37229 12624 37315
rect 6049 37087 6125 37173
rect 10425 37200 11495 37210
rect 10425 37144 10435 37200
rect 10491 37144 10577 37200
rect 10633 37144 10719 37200
rect 10775 37144 10861 37200
rect 10917 37144 11003 37200
rect 11059 37144 11145 37200
rect 11201 37144 11287 37200
rect 11343 37144 11429 37200
rect 11485 37144 11495 37200
rect 10425 37134 11495 37144
rect 12406 37173 12416 37229
rect 12472 37173 12558 37229
rect 12614 37173 12624 37229
rect 6049 37031 6059 37087
rect 6115 37031 6125 37087
rect 6049 36945 6125 37031
rect 6049 36889 6059 36945
rect 6115 36889 6125 36945
rect 6049 36803 6125 36889
rect 6049 36747 6059 36803
rect 6115 36747 6125 36803
rect 6049 36661 6125 36747
rect 6049 36605 6059 36661
rect 6115 36605 6125 36661
rect 6049 36519 6125 36605
rect 6049 36463 6059 36519
rect 6115 36463 6125 36519
rect 6049 36453 6125 36463
rect 12406 37087 12624 37173
rect 12406 37031 12416 37087
rect 12472 37031 12558 37087
rect 12614 37031 12624 37087
rect 12406 36945 12624 37031
rect 12406 36889 12416 36945
rect 12472 36889 12558 36945
rect 12614 36889 12624 36945
rect 12406 36803 12624 36889
rect 12406 36747 12416 36803
rect 12472 36747 12558 36803
rect 12614 36747 12624 36803
rect 12406 36661 12624 36747
rect 12406 36605 12416 36661
rect 12472 36605 12558 36661
rect 12614 36605 12624 36661
rect 12406 36519 12624 36605
rect 12406 36463 12416 36519
rect 12472 36463 12558 36519
rect 12614 36463 12624 36519
rect 12406 36453 12624 36463
rect 14942 37797 15018 37807
rect 14942 37741 14952 37797
rect 15008 37741 15018 37797
rect 14942 37655 15018 37741
rect 14942 37599 14952 37655
rect 15008 37599 15018 37655
rect 14942 37513 15018 37599
rect 14942 37457 14952 37513
rect 15008 37457 15018 37513
rect 14942 37371 15018 37457
rect 14942 37315 14952 37371
rect 15008 37315 15018 37371
rect 14942 37229 15018 37315
rect 14942 37173 14952 37229
rect 15008 37173 15018 37229
rect 14942 37087 15018 37173
rect 14942 37031 14952 37087
rect 15008 37031 15018 37087
rect 14942 36945 15018 37031
rect 14942 36889 14952 36945
rect 15008 36889 15018 36945
rect 14942 36803 15018 36889
rect 14942 36747 14952 36803
rect 15008 36747 15018 36803
rect 14942 36661 15018 36747
rect 14942 36605 14952 36661
rect 15008 36605 15018 36661
rect 14942 36519 15018 36605
rect 14942 36463 14952 36519
rect 15008 36463 15018 36519
rect 14942 36453 15018 36463
rect 165 36178 383 36188
rect 165 36122 175 36178
rect 231 36122 317 36178
rect 373 36122 383 36178
rect 165 36036 383 36122
rect 165 35980 175 36036
rect 231 35980 317 36036
rect 373 35980 383 36036
rect 165 35894 383 35980
rect 165 35838 175 35894
rect 231 35838 317 35894
rect 373 35838 383 35894
rect 165 35752 383 35838
rect 165 35696 175 35752
rect 231 35696 317 35752
rect 373 35696 383 35752
rect 165 35610 383 35696
rect 3990 35716 4066 35726
rect 3990 35660 4000 35716
rect 4056 35660 4066 35716
rect 165 35554 175 35610
rect 231 35554 317 35610
rect 373 35554 383 35610
rect 165 35468 383 35554
rect 165 35412 175 35468
rect 231 35412 317 35468
rect 373 35412 383 35468
rect 165 35326 383 35412
rect 165 35270 175 35326
rect 231 35270 317 35326
rect 373 35270 383 35326
rect 165 35184 383 35270
rect 165 35128 175 35184
rect 231 35128 317 35184
rect 373 35128 383 35184
rect 165 35042 383 35128
rect 165 34986 175 35042
rect 231 34986 317 35042
rect 373 34986 383 35042
rect 165 34900 383 34986
rect 165 34844 175 34900
rect 231 34844 317 34900
rect 373 34844 383 34900
rect 165 34758 383 34844
rect 165 34702 175 34758
rect 231 34702 317 34758
rect 373 34702 383 34758
rect 165 34616 383 34702
rect 165 34560 175 34616
rect 231 34560 317 34616
rect 373 34560 383 34616
rect 165 34474 383 34560
rect 165 34418 175 34474
rect 231 34418 317 34474
rect 373 34418 383 34474
rect 165 34332 383 34418
rect 165 34276 175 34332
rect 231 34276 317 34332
rect 373 34276 383 34332
rect 165 34190 383 34276
rect 165 34134 175 34190
rect 231 34134 317 34190
rect 373 34134 383 34190
rect 165 34048 383 34134
rect 165 33992 175 34048
rect 231 33992 317 34048
rect 373 33992 383 34048
rect 165 33906 383 33992
rect 165 33850 175 33906
rect 231 33850 317 33906
rect 373 33850 383 33906
rect 165 33764 383 33850
rect 165 33708 175 33764
rect 231 33708 317 33764
rect 373 33708 383 33764
rect 165 33622 383 33708
rect 486 35617 562 35627
rect 486 35561 496 35617
rect 552 35561 562 35617
rect 486 35475 562 35561
rect 486 35419 496 35475
rect 552 35419 562 35475
rect 486 35333 562 35419
rect 486 35277 496 35333
rect 552 35277 562 35333
rect 486 35191 562 35277
rect 486 35135 496 35191
rect 552 35135 562 35191
rect 486 35049 562 35135
rect 486 34993 496 35049
rect 552 34993 562 35049
rect 486 34907 562 34993
rect 486 34851 496 34907
rect 552 34851 562 34907
rect 486 34765 562 34851
rect 486 34709 496 34765
rect 552 34709 562 34765
rect 486 34623 562 34709
rect 486 34567 496 34623
rect 552 34567 562 34623
rect 486 34481 562 34567
rect 486 34425 496 34481
rect 552 34425 562 34481
rect 486 34339 562 34425
rect 486 34283 496 34339
rect 552 34283 562 34339
rect 486 34197 562 34283
rect 486 34141 496 34197
rect 552 34141 562 34197
rect 486 34055 562 34141
rect 724 35612 800 35622
rect 724 35556 734 35612
rect 790 35556 800 35612
rect 724 35470 800 35556
rect 724 35414 734 35470
rect 790 35414 800 35470
rect 724 35328 800 35414
rect 724 35272 734 35328
rect 790 35272 800 35328
rect 724 35186 800 35272
rect 724 35130 734 35186
rect 790 35130 800 35186
rect 724 35044 800 35130
rect 724 34988 734 35044
rect 790 34988 800 35044
rect 724 34902 800 34988
rect 724 34846 734 34902
rect 790 34846 800 34902
rect 724 34760 800 34846
rect 724 34704 734 34760
rect 790 34704 800 34760
rect 724 34618 800 34704
rect 724 34562 734 34618
rect 790 34562 800 34618
rect 724 34476 800 34562
rect 724 34420 734 34476
rect 790 34420 800 34476
rect 724 34334 800 34420
rect 724 34278 734 34334
rect 790 34278 800 34334
rect 724 34192 800 34278
rect 724 34136 734 34192
rect 790 34136 800 34192
rect 724 34126 800 34136
rect 3092 35612 3168 35622
rect 3092 35556 3102 35612
rect 3158 35556 3168 35612
rect 3092 35470 3168 35556
rect 3092 35414 3102 35470
rect 3158 35414 3168 35470
rect 3092 35328 3168 35414
rect 3092 35272 3102 35328
rect 3158 35272 3168 35328
rect 3092 35186 3168 35272
rect 3092 35130 3102 35186
rect 3158 35130 3168 35186
rect 3092 35044 3168 35130
rect 3092 34988 3102 35044
rect 3158 34988 3168 35044
rect 3092 34902 3168 34988
rect 3092 34846 3102 34902
rect 3158 34846 3168 34902
rect 3092 34760 3168 34846
rect 3092 34704 3102 34760
rect 3158 34704 3168 34760
rect 3092 34618 3168 34704
rect 3092 34562 3102 34618
rect 3158 34562 3168 34618
rect 3092 34476 3168 34562
rect 3092 34420 3102 34476
rect 3158 34420 3168 34476
rect 3092 34334 3168 34420
rect 3092 34278 3102 34334
rect 3158 34278 3168 34334
rect 3092 34192 3168 34278
rect 3092 34136 3102 34192
rect 3158 34136 3168 34192
rect 3092 34126 3168 34136
rect 3990 35574 4066 35660
rect 10998 35716 11074 35726
rect 10998 35660 11008 35716
rect 11064 35660 11074 35716
rect 3990 35518 4000 35574
rect 4056 35518 4066 35574
rect 3990 35432 4066 35518
rect 3990 35376 4000 35432
rect 4056 35376 4066 35432
rect 3990 35290 4066 35376
rect 3990 35234 4000 35290
rect 4056 35234 4066 35290
rect 3990 35148 4066 35234
rect 3990 35092 4000 35148
rect 4056 35092 4066 35148
rect 3990 35006 4066 35092
rect 3990 34950 4000 35006
rect 4056 34950 4066 35006
rect 3990 34864 4066 34950
rect 3990 34808 4000 34864
rect 4056 34808 4066 34864
rect 3990 34722 4066 34808
rect 3990 34666 4000 34722
rect 4056 34666 4066 34722
rect 3990 34580 4066 34666
rect 3990 34524 4000 34580
rect 4056 34524 4066 34580
rect 3990 34438 4066 34524
rect 3990 34382 4000 34438
rect 4056 34382 4066 34438
rect 3990 34296 4066 34382
rect 3990 34240 4000 34296
rect 4056 34240 4066 34296
rect 3990 34154 4066 34240
rect 486 33999 496 34055
rect 552 33999 562 34055
rect 486 33913 562 33999
rect 486 33857 496 33913
rect 552 33857 562 33913
rect 486 33771 562 33857
rect 486 33715 496 33771
rect 552 33715 562 33771
rect 486 33705 562 33715
rect 3990 34098 4000 34154
rect 4056 34098 4066 34154
rect 4888 35612 4964 35622
rect 4888 35556 4898 35612
rect 4954 35556 4964 35612
rect 4888 35470 4964 35556
rect 4888 35414 4898 35470
rect 4954 35414 4964 35470
rect 4888 35328 4964 35414
rect 4888 35272 4898 35328
rect 4954 35272 4964 35328
rect 4888 35186 4964 35272
rect 4888 35130 4898 35186
rect 4954 35130 4964 35186
rect 4888 35044 4964 35130
rect 4888 34988 4898 35044
rect 4954 34988 4964 35044
rect 4888 34902 4964 34988
rect 4888 34846 4898 34902
rect 4954 34846 4964 34902
rect 4888 34760 4964 34846
rect 4888 34704 4898 34760
rect 4954 34704 4964 34760
rect 4888 34618 4964 34704
rect 4888 34562 4898 34618
rect 4954 34562 4964 34618
rect 4888 34476 4964 34562
rect 4888 34420 4898 34476
rect 4954 34420 4964 34476
rect 4888 34334 4964 34420
rect 4888 34278 4898 34334
rect 4954 34278 4964 34334
rect 4888 34192 4964 34278
rect 4888 34136 4898 34192
rect 4954 34136 4964 34192
rect 4888 34126 4964 34136
rect 8671 35612 8747 35622
rect 8671 35556 8681 35612
rect 8737 35556 8747 35612
rect 8671 35470 8747 35556
rect 8671 35414 8681 35470
rect 8737 35414 8747 35470
rect 8671 35328 8747 35414
rect 8671 35272 8681 35328
rect 8737 35272 8747 35328
rect 8671 35186 8747 35272
rect 8671 35130 8681 35186
rect 8737 35130 8747 35186
rect 8671 35044 8747 35130
rect 8671 34988 8681 35044
rect 8737 34988 8747 35044
rect 8671 34902 8747 34988
rect 8671 34846 8681 34902
rect 8737 34846 8747 34902
rect 8671 34760 8747 34846
rect 8671 34704 8681 34760
rect 8737 34704 8747 34760
rect 8671 34618 8747 34704
rect 8671 34562 8681 34618
rect 8737 34562 8747 34618
rect 8671 34476 8747 34562
rect 8671 34420 8681 34476
rect 8737 34420 8747 34476
rect 8671 34334 8747 34420
rect 8671 34278 8681 34334
rect 8737 34278 8747 34334
rect 8671 34192 8747 34278
rect 8671 34136 8681 34192
rect 8737 34136 8747 34192
rect 8671 34126 8747 34136
rect 10100 35612 10176 35622
rect 10100 35556 10110 35612
rect 10166 35556 10176 35612
rect 10100 35470 10176 35556
rect 10100 35414 10110 35470
rect 10166 35414 10176 35470
rect 10100 35328 10176 35414
rect 10100 35272 10110 35328
rect 10166 35272 10176 35328
rect 10100 35186 10176 35272
rect 10100 35130 10110 35186
rect 10166 35130 10176 35186
rect 10100 35044 10176 35130
rect 10100 34988 10110 35044
rect 10166 34988 10176 35044
rect 10100 34902 10176 34988
rect 10100 34846 10110 34902
rect 10166 34846 10176 34902
rect 10100 34760 10176 34846
rect 10100 34704 10110 34760
rect 10166 34704 10176 34760
rect 10100 34618 10176 34704
rect 10100 34562 10110 34618
rect 10166 34562 10176 34618
rect 10100 34476 10176 34562
rect 10100 34420 10110 34476
rect 10166 34420 10176 34476
rect 10100 34334 10176 34420
rect 10100 34278 10110 34334
rect 10166 34278 10176 34334
rect 10100 34192 10176 34278
rect 10100 34136 10110 34192
rect 10166 34136 10176 34192
rect 10100 34126 10176 34136
rect 10998 35574 11074 35660
rect 10998 35518 11008 35574
rect 11064 35518 11074 35574
rect 10998 35432 11074 35518
rect 10998 35376 11008 35432
rect 11064 35376 11074 35432
rect 10998 35290 11074 35376
rect 10998 35234 11008 35290
rect 11064 35234 11074 35290
rect 10998 35148 11074 35234
rect 10998 35092 11008 35148
rect 11064 35092 11074 35148
rect 10998 35006 11074 35092
rect 10998 34950 11008 35006
rect 11064 34950 11074 35006
rect 10998 34864 11074 34950
rect 10998 34808 11008 34864
rect 11064 34808 11074 34864
rect 10998 34722 11074 34808
rect 10998 34666 11008 34722
rect 11064 34666 11074 34722
rect 10998 34580 11074 34666
rect 10998 34524 11008 34580
rect 11064 34524 11074 34580
rect 10998 34438 11074 34524
rect 10998 34382 11008 34438
rect 11064 34382 11074 34438
rect 10998 34296 11074 34382
rect 10998 34240 11008 34296
rect 11064 34240 11074 34296
rect 10998 34154 11074 34240
rect 3990 34012 4066 34098
rect 3990 33956 4000 34012
rect 4056 33956 4066 34012
rect 3990 33870 4066 33956
rect 3990 33814 4000 33870
rect 4056 33814 4066 33870
rect 3990 33728 4066 33814
rect 165 33566 175 33622
rect 231 33566 317 33622
rect 373 33566 383 33622
rect 165 33480 383 33566
rect 165 33424 175 33480
rect 231 33424 317 33480
rect 373 33424 383 33480
rect 165 33338 383 33424
rect 165 33282 175 33338
rect 231 33282 317 33338
rect 373 33282 383 33338
rect 165 33272 383 33282
rect 3990 33672 4000 33728
rect 4056 33672 4066 33728
rect 3990 33586 4066 33672
rect 3990 33530 4000 33586
rect 4056 33530 4066 33586
rect 3990 33444 4066 33530
rect 3990 33388 4000 33444
rect 4056 33388 4066 33444
rect 3990 33302 4066 33388
rect 3990 33246 4000 33302
rect 4056 33246 4066 33302
rect 3990 33236 4066 33246
rect 10998 34098 11008 34154
rect 11064 34098 11074 34154
rect 11896 35612 11972 35622
rect 11896 35556 11906 35612
rect 11962 35556 11972 35612
rect 11896 35470 11972 35556
rect 11896 35414 11906 35470
rect 11962 35414 11972 35470
rect 11896 35328 11972 35414
rect 11896 35272 11906 35328
rect 11962 35272 11972 35328
rect 11896 35186 11972 35272
rect 11896 35130 11906 35186
rect 11962 35130 11972 35186
rect 11896 35044 11972 35130
rect 11896 34988 11906 35044
rect 11962 34988 11972 35044
rect 11896 34902 11972 34988
rect 11896 34846 11906 34902
rect 11962 34846 11972 34902
rect 11896 34760 11972 34846
rect 11896 34704 11906 34760
rect 11962 34704 11972 34760
rect 11896 34618 11972 34704
rect 11896 34562 11906 34618
rect 11962 34562 11972 34618
rect 11896 34476 11972 34562
rect 11896 34420 11906 34476
rect 11962 34420 11972 34476
rect 11896 34334 11972 34420
rect 11896 34278 11906 34334
rect 11962 34278 11972 34334
rect 11896 34192 11972 34278
rect 11896 34136 11906 34192
rect 11962 34136 11972 34192
rect 11896 34126 11972 34136
rect 10998 34012 11074 34098
rect 10998 33956 11008 34012
rect 11064 33956 11074 34012
rect 10998 33870 11074 33956
rect 10998 33814 11008 33870
rect 11064 33814 11074 33870
rect 10998 33728 11074 33814
rect 10998 33672 11008 33728
rect 11064 33672 11074 33728
rect 10998 33586 11074 33672
rect 10998 33530 11008 33586
rect 11064 33530 11074 33586
rect 10998 33444 11074 33530
rect 10998 33388 11008 33444
rect 11064 33388 11074 33444
rect 10998 33302 11074 33388
rect 10998 33246 11008 33302
rect 11064 33246 11074 33302
rect 10998 33236 11074 33246
rect 486 32978 562 32988
rect 486 32922 496 32978
rect 552 32922 562 32978
rect 486 32836 562 32922
rect 486 32780 496 32836
rect 552 32780 562 32836
rect 486 32694 562 32780
rect 486 32638 496 32694
rect 552 32638 562 32694
rect 486 32552 562 32638
rect 486 32496 496 32552
rect 552 32496 562 32552
rect 14400 32978 14760 32988
rect 14400 32922 14410 32978
rect 14466 32922 14552 32978
rect 14608 32922 14694 32978
rect 14750 32922 14760 32978
rect 14400 32836 14760 32922
rect 14400 32780 14410 32836
rect 14466 32780 14552 32836
rect 14608 32780 14694 32836
rect 14750 32780 14760 32836
rect 14400 32694 14760 32780
rect 14400 32638 14410 32694
rect 14466 32638 14552 32694
rect 14608 32638 14694 32694
rect 14750 32638 14760 32694
rect 14400 32552 14760 32638
rect 486 32410 562 32496
rect 486 32354 496 32410
rect 552 32354 562 32410
rect 486 32268 562 32354
rect 3990 32535 4066 32545
rect 3990 32479 4000 32535
rect 4056 32479 4066 32535
rect 3990 32393 4066 32479
rect 3990 32337 4000 32393
rect 4056 32337 4066 32393
rect 486 32212 496 32268
rect 552 32212 562 32268
rect 486 32126 562 32212
rect 486 32070 496 32126
rect 552 32070 562 32126
rect 486 31984 562 32070
rect 486 31928 496 31984
rect 552 31928 562 31984
rect 486 31842 562 31928
rect 486 31786 496 31842
rect 552 31786 562 31842
rect 486 31700 562 31786
rect 486 31644 496 31700
rect 552 31644 562 31700
rect 486 31558 562 31644
rect 486 31502 496 31558
rect 552 31502 562 31558
rect 486 31416 562 31502
rect 486 31360 496 31416
rect 552 31360 562 31416
rect 486 31274 562 31360
rect 486 31218 496 31274
rect 552 31218 562 31274
rect 486 31132 562 31218
rect 486 31076 496 31132
rect 552 31076 562 31132
rect 486 30990 562 31076
rect 486 30934 496 30990
rect 552 30934 562 30990
rect 486 30848 562 30934
rect 486 30792 496 30848
rect 552 30792 562 30848
rect 486 30706 562 30792
rect 486 30650 496 30706
rect 552 30650 562 30706
rect 486 30564 562 30650
rect 486 30508 496 30564
rect 552 30508 562 30564
rect 486 30422 562 30508
rect 486 30366 496 30422
rect 552 30366 562 30422
rect 486 30280 562 30366
rect 486 30224 496 30280
rect 552 30224 562 30280
rect 486 30138 562 30224
rect 486 30082 496 30138
rect 552 30082 562 30138
rect 968 32322 1044 32332
rect 968 32266 978 32322
rect 1034 32266 1044 32322
rect 968 32180 1044 32266
rect 968 32124 978 32180
rect 1034 32124 1044 32180
rect 968 32038 1044 32124
rect 968 31982 978 32038
rect 1034 31982 1044 32038
rect 968 31896 1044 31982
rect 968 31840 978 31896
rect 1034 31840 1044 31896
rect 968 31754 1044 31840
rect 968 31698 978 31754
rect 1034 31698 1044 31754
rect 968 31612 1044 31698
rect 968 31556 978 31612
rect 1034 31556 1044 31612
rect 968 31470 1044 31556
rect 968 31414 978 31470
rect 1034 31414 1044 31470
rect 968 31328 1044 31414
rect 968 31272 978 31328
rect 1034 31272 1044 31328
rect 968 31186 1044 31272
rect 968 31130 978 31186
rect 1034 31130 1044 31186
rect 968 31044 1044 31130
rect 968 30988 978 31044
rect 1034 30988 1044 31044
rect 968 30902 1044 30988
rect 968 30846 978 30902
rect 1034 30846 1044 30902
rect 968 30760 1044 30846
rect 968 30704 978 30760
rect 1034 30704 1044 30760
rect 968 30618 1044 30704
rect 968 30562 978 30618
rect 1034 30562 1044 30618
rect 968 30476 1044 30562
rect 968 30420 978 30476
rect 1034 30420 1044 30476
rect 968 30334 1044 30420
rect 968 30278 978 30334
rect 1034 30278 1044 30334
rect 968 30192 1044 30278
rect 968 30136 978 30192
rect 1034 30136 1044 30192
rect 968 30126 1044 30136
rect 2360 32322 2436 32332
rect 2360 32266 2370 32322
rect 2426 32266 2436 32322
rect 2360 32180 2436 32266
rect 2360 32124 2370 32180
rect 2426 32124 2436 32180
rect 2360 32038 2436 32124
rect 2360 31982 2370 32038
rect 2426 31982 2436 32038
rect 2360 31896 2436 31982
rect 2360 31840 2370 31896
rect 2426 31840 2436 31896
rect 2360 31754 2436 31840
rect 2360 31698 2370 31754
rect 2426 31698 2436 31754
rect 2360 31612 2436 31698
rect 2360 31556 2370 31612
rect 2426 31556 2436 31612
rect 2360 31470 2436 31556
rect 2360 31414 2370 31470
rect 2426 31414 2436 31470
rect 2360 31328 2436 31414
rect 2360 31272 2370 31328
rect 2426 31272 2436 31328
rect 2360 31186 2436 31272
rect 2360 31130 2370 31186
rect 2426 31130 2436 31186
rect 2360 31044 2436 31130
rect 2360 30988 2370 31044
rect 2426 30988 2436 31044
rect 2360 30902 2436 30988
rect 2360 30846 2370 30902
rect 2426 30846 2436 30902
rect 2360 30760 2436 30846
rect 2360 30704 2370 30760
rect 2426 30704 2436 30760
rect 2360 30618 2436 30704
rect 2360 30562 2370 30618
rect 2426 30562 2436 30618
rect 2360 30476 2436 30562
rect 2360 30420 2370 30476
rect 2426 30420 2436 30476
rect 2360 30334 2436 30420
rect 2360 30278 2370 30334
rect 2426 30278 2436 30334
rect 2360 30192 2436 30278
rect 2360 30136 2370 30192
rect 2426 30136 2436 30192
rect 2360 30126 2436 30136
rect 2776 32322 2852 32332
rect 2776 32266 2786 32322
rect 2842 32266 2852 32322
rect 2776 32180 2852 32266
rect 2776 32124 2786 32180
rect 2842 32124 2852 32180
rect 2776 32038 2852 32124
rect 2776 31982 2786 32038
rect 2842 31982 2852 32038
rect 2776 31896 2852 31982
rect 2776 31840 2786 31896
rect 2842 31840 2852 31896
rect 2776 31754 2852 31840
rect 2776 31698 2786 31754
rect 2842 31698 2852 31754
rect 2776 31612 2852 31698
rect 2776 31556 2786 31612
rect 2842 31556 2852 31612
rect 2776 31470 2852 31556
rect 2776 31414 2786 31470
rect 2842 31414 2852 31470
rect 2776 31328 2852 31414
rect 2776 31272 2786 31328
rect 2842 31272 2852 31328
rect 2776 31186 2852 31272
rect 2776 31130 2786 31186
rect 2842 31130 2852 31186
rect 2776 31044 2852 31130
rect 2776 30988 2786 31044
rect 2842 30988 2852 31044
rect 2776 30902 2852 30988
rect 2776 30846 2786 30902
rect 2842 30846 2852 30902
rect 2776 30760 2852 30846
rect 2776 30704 2786 30760
rect 2842 30704 2852 30760
rect 2776 30618 2852 30704
rect 3264 32323 3340 32333
rect 3264 32267 3274 32323
rect 3330 32267 3340 32323
rect 3264 32181 3340 32267
rect 3264 32125 3274 32181
rect 3330 32125 3340 32181
rect 3264 32039 3340 32125
rect 3264 31983 3274 32039
rect 3330 31983 3340 32039
rect 3264 31897 3340 31983
rect 3264 31841 3274 31897
rect 3330 31841 3340 31897
rect 3264 31755 3340 31841
rect 3264 31699 3274 31755
rect 3330 31699 3340 31755
rect 3264 31613 3340 31699
rect 3264 31557 3274 31613
rect 3330 31557 3340 31613
rect 3264 31471 3340 31557
rect 3264 31415 3274 31471
rect 3330 31415 3340 31471
rect 3264 31329 3340 31415
rect 3264 31273 3274 31329
rect 3330 31273 3340 31329
rect 3264 31187 3340 31273
rect 3264 31131 3274 31187
rect 3330 31131 3340 31187
rect 3264 31045 3340 31131
rect 3264 30989 3274 31045
rect 3330 30989 3340 31045
rect 3264 30903 3340 30989
rect 3264 30847 3274 30903
rect 3330 30847 3340 30903
rect 3264 30761 3340 30847
rect 3264 30705 3274 30761
rect 3330 30705 3340 30761
rect 3264 30695 3340 30705
rect 3752 32272 3828 32282
rect 3752 32216 3762 32272
rect 3818 32216 3828 32272
rect 3752 32130 3828 32216
rect 3752 32074 3762 32130
rect 3818 32074 3828 32130
rect 3752 31988 3828 32074
rect 3752 31932 3762 31988
rect 3818 31932 3828 31988
rect 3752 31846 3828 31932
rect 3752 31790 3762 31846
rect 3818 31790 3828 31846
rect 3752 31704 3828 31790
rect 3752 31648 3762 31704
rect 3818 31648 3828 31704
rect 3752 31562 3828 31648
rect 3752 31506 3762 31562
rect 3818 31506 3828 31562
rect 3752 31420 3828 31506
rect 3752 31364 3762 31420
rect 3818 31364 3828 31420
rect 3752 31278 3828 31364
rect 3752 31222 3762 31278
rect 3818 31222 3828 31278
rect 3752 31136 3828 31222
rect 3752 31080 3762 31136
rect 3818 31080 3828 31136
rect 3752 30994 3828 31080
rect 3752 30938 3762 30994
rect 3818 30938 3828 30994
rect 3752 30852 3828 30938
rect 3752 30796 3762 30852
rect 3818 30796 3828 30852
rect 3752 30710 3828 30796
rect 3752 30654 3762 30710
rect 3818 30654 3828 30710
rect 3752 30644 3828 30654
rect 3990 32251 4066 32337
rect 10998 32535 11074 32545
rect 10998 32479 11008 32535
rect 11064 32479 11074 32535
rect 10998 32393 11074 32479
rect 10998 32337 11008 32393
rect 11064 32337 11074 32393
rect 4716 32323 4792 32333
rect 3990 32195 4000 32251
rect 4056 32195 4066 32251
rect 3990 32109 4066 32195
rect 3990 32053 4000 32109
rect 4056 32053 4066 32109
rect 3990 31967 4066 32053
rect 3990 31911 4000 31967
rect 4056 31911 4066 31967
rect 3990 31825 4066 31911
rect 3990 31769 4000 31825
rect 4056 31769 4066 31825
rect 3990 31683 4066 31769
rect 3990 31627 4000 31683
rect 4056 31627 4066 31683
rect 3990 31541 4066 31627
rect 3990 31485 4000 31541
rect 4056 31485 4066 31541
rect 3990 31399 4066 31485
rect 3990 31343 4000 31399
rect 4056 31343 4066 31399
rect 3990 31257 4066 31343
rect 3990 31201 4000 31257
rect 4056 31201 4066 31257
rect 3990 31115 4066 31201
rect 3990 31059 4000 31115
rect 4056 31059 4066 31115
rect 3990 30973 4066 31059
rect 3990 30917 4000 30973
rect 4056 30917 4066 30973
rect 3990 30831 4066 30917
rect 3990 30775 4000 30831
rect 4056 30775 4066 30831
rect 3990 30689 4066 30775
rect 3990 30633 4000 30689
rect 4056 30633 4066 30689
rect 4228 32272 4304 32282
rect 4228 32216 4238 32272
rect 4294 32216 4304 32272
rect 4228 32130 4304 32216
rect 4228 32074 4238 32130
rect 4294 32074 4304 32130
rect 4228 31988 4304 32074
rect 4228 31932 4238 31988
rect 4294 31932 4304 31988
rect 4228 31846 4304 31932
rect 4228 31790 4238 31846
rect 4294 31790 4304 31846
rect 4228 31704 4304 31790
rect 4228 31648 4238 31704
rect 4294 31648 4304 31704
rect 4228 31562 4304 31648
rect 4228 31506 4238 31562
rect 4294 31506 4304 31562
rect 4228 31420 4304 31506
rect 4228 31364 4238 31420
rect 4294 31364 4304 31420
rect 4228 31278 4304 31364
rect 4228 31222 4238 31278
rect 4294 31222 4304 31278
rect 4228 31136 4304 31222
rect 4228 31080 4238 31136
rect 4294 31080 4304 31136
rect 4228 30994 4304 31080
rect 4228 30938 4238 30994
rect 4294 30938 4304 30994
rect 4228 30852 4304 30938
rect 4228 30796 4238 30852
rect 4294 30796 4304 30852
rect 4228 30710 4304 30796
rect 4228 30654 4238 30710
rect 4294 30654 4304 30710
rect 4716 32267 4726 32323
rect 4782 32267 4792 32323
rect 4716 32181 4792 32267
rect 4716 32125 4726 32181
rect 4782 32125 4792 32181
rect 4716 32039 4792 32125
rect 4716 31983 4726 32039
rect 4782 31983 4792 32039
rect 4716 31897 4792 31983
rect 4716 31841 4726 31897
rect 4782 31841 4792 31897
rect 4716 31755 4792 31841
rect 4716 31699 4726 31755
rect 4782 31699 4792 31755
rect 4716 31613 4792 31699
rect 4716 31557 4726 31613
rect 4782 31557 4792 31613
rect 4716 31471 4792 31557
rect 4716 31415 4726 31471
rect 4782 31415 4792 31471
rect 4716 31329 4792 31415
rect 4716 31273 4726 31329
rect 4782 31273 4792 31329
rect 4716 31187 4792 31273
rect 4716 31131 4726 31187
rect 4782 31131 4792 31187
rect 4716 31045 4792 31131
rect 4716 30989 4726 31045
rect 4782 30989 4792 31045
rect 4716 30903 4792 30989
rect 4716 30847 4726 30903
rect 4782 30847 4792 30903
rect 4716 30761 4792 30847
rect 4716 30705 4726 30761
rect 4782 30705 4792 30761
rect 4716 30695 4792 30705
rect 5204 32323 5280 32333
rect 5204 32267 5214 32323
rect 5270 32267 5280 32323
rect 5204 32181 5280 32267
rect 5204 32125 5214 32181
rect 5270 32125 5280 32181
rect 5204 32039 5280 32125
rect 5204 31983 5214 32039
rect 5270 31983 5280 32039
rect 5204 31897 5280 31983
rect 5204 31841 5214 31897
rect 5270 31841 5280 31897
rect 5204 31755 5280 31841
rect 5204 31699 5214 31755
rect 5270 31699 5280 31755
rect 5204 31613 5280 31699
rect 5204 31557 5214 31613
rect 5270 31557 5280 31613
rect 5204 31471 5280 31557
rect 5204 31415 5214 31471
rect 5270 31415 5280 31471
rect 5204 31329 5280 31415
rect 5204 31273 5214 31329
rect 5270 31273 5280 31329
rect 5204 31187 5280 31273
rect 5204 31131 5214 31187
rect 5270 31131 5280 31187
rect 5204 31045 5280 31131
rect 5204 30989 5214 31045
rect 5270 30989 5280 31045
rect 5204 30903 5280 30989
rect 5204 30847 5214 30903
rect 5270 30847 5280 30903
rect 5204 30761 5280 30847
rect 5204 30705 5214 30761
rect 5270 30705 5280 30761
rect 5204 30695 5280 30705
rect 5620 32323 5696 32333
rect 5620 32267 5630 32323
rect 5686 32267 5696 32323
rect 5620 32181 5696 32267
rect 5620 32125 5630 32181
rect 5686 32125 5696 32181
rect 5620 32039 5696 32125
rect 5620 31983 5630 32039
rect 5686 31983 5696 32039
rect 5620 31897 5696 31983
rect 5620 31841 5630 31897
rect 5686 31841 5696 31897
rect 5620 31755 5696 31841
rect 5620 31699 5630 31755
rect 5686 31699 5696 31755
rect 5620 31613 5696 31699
rect 5620 31557 5630 31613
rect 5686 31557 5696 31613
rect 5620 31471 5696 31557
rect 5620 31415 5630 31471
rect 5686 31415 5696 31471
rect 5620 31329 5696 31415
rect 5620 31273 5630 31329
rect 5686 31273 5696 31329
rect 5620 31187 5696 31273
rect 5620 31131 5630 31187
rect 5686 31131 5696 31187
rect 5620 31045 5696 31131
rect 5620 30989 5630 31045
rect 5686 30989 5696 31045
rect 5620 30903 5696 30989
rect 5620 30847 5630 30903
rect 5686 30847 5696 30903
rect 5620 30761 5696 30847
rect 5620 30705 5630 30761
rect 5686 30705 5696 30761
rect 5620 30695 5696 30705
rect 7012 32322 7088 32332
rect 7012 32266 7022 32322
rect 7078 32266 7088 32322
rect 7012 32180 7088 32266
rect 7012 32124 7022 32180
rect 7078 32124 7088 32180
rect 7012 32038 7088 32124
rect 7012 31982 7022 32038
rect 7078 31982 7088 32038
rect 7012 31896 7088 31982
rect 7012 31840 7022 31896
rect 7078 31840 7088 31896
rect 7012 31754 7088 31840
rect 7012 31698 7022 31754
rect 7078 31698 7088 31754
rect 7012 31612 7088 31698
rect 7012 31556 7022 31612
rect 7078 31556 7088 31612
rect 7012 31470 7088 31556
rect 7012 31414 7022 31470
rect 7078 31414 7088 31470
rect 7012 31328 7088 31414
rect 7012 31272 7022 31328
rect 7078 31272 7088 31328
rect 7012 31186 7088 31272
rect 7012 31130 7022 31186
rect 7078 31130 7088 31186
rect 7012 31044 7088 31130
rect 7012 30988 7022 31044
rect 7078 30988 7088 31044
rect 7012 30902 7088 30988
rect 7012 30846 7022 30902
rect 7078 30846 7088 30902
rect 7012 30760 7088 30846
rect 7012 30704 7022 30760
rect 7078 30704 7088 30760
rect 4228 30644 4304 30654
rect 3990 30623 4066 30633
rect 2776 30562 2786 30618
rect 2842 30562 2852 30618
rect 2776 30476 2852 30562
rect 2776 30420 2786 30476
rect 2842 30420 2852 30476
rect 2776 30334 2852 30420
rect 2776 30278 2786 30334
rect 2842 30278 2852 30334
rect 2776 30192 2852 30278
rect 2776 30136 2786 30192
rect 2842 30136 2852 30192
rect 2776 30126 2852 30136
rect 7012 30618 7088 30704
rect 7012 30562 7022 30618
rect 7078 30562 7088 30618
rect 7012 30476 7088 30562
rect 7012 30420 7022 30476
rect 7078 30420 7088 30476
rect 7012 30334 7088 30420
rect 7012 30278 7022 30334
rect 7078 30278 7088 30334
rect 7012 30192 7088 30278
rect 7012 30136 7022 30192
rect 7078 30136 7088 30192
rect 7012 30126 7088 30136
rect 7976 32322 8052 32332
rect 7976 32266 7986 32322
rect 8042 32266 8052 32322
rect 7976 32180 8052 32266
rect 7976 32124 7986 32180
rect 8042 32124 8052 32180
rect 7976 32038 8052 32124
rect 7976 31982 7986 32038
rect 8042 31982 8052 32038
rect 7976 31896 8052 31982
rect 7976 31840 7986 31896
rect 8042 31840 8052 31896
rect 7976 31754 8052 31840
rect 7976 31698 7986 31754
rect 8042 31698 8052 31754
rect 7976 31612 8052 31698
rect 7976 31556 7986 31612
rect 8042 31556 8052 31612
rect 7976 31470 8052 31556
rect 7976 31414 7986 31470
rect 8042 31414 8052 31470
rect 7976 31328 8052 31414
rect 7976 31272 7986 31328
rect 8042 31272 8052 31328
rect 7976 31186 8052 31272
rect 7976 31130 7986 31186
rect 8042 31130 8052 31186
rect 7976 31044 8052 31130
rect 7976 30988 7986 31044
rect 8042 30988 8052 31044
rect 7976 30902 8052 30988
rect 7976 30846 7986 30902
rect 8042 30846 8052 30902
rect 7976 30760 8052 30846
rect 7976 30704 7986 30760
rect 8042 30704 8052 30760
rect 7976 30618 8052 30704
rect 9368 32323 9444 32333
rect 9368 32267 9378 32323
rect 9434 32267 9444 32323
rect 9368 32181 9444 32267
rect 9368 32125 9378 32181
rect 9434 32125 9444 32181
rect 9368 32039 9444 32125
rect 9368 31983 9378 32039
rect 9434 31983 9444 32039
rect 9368 31897 9444 31983
rect 9368 31841 9378 31897
rect 9434 31841 9444 31897
rect 9368 31755 9444 31841
rect 9368 31699 9378 31755
rect 9434 31699 9444 31755
rect 9368 31613 9444 31699
rect 9368 31557 9378 31613
rect 9434 31557 9444 31613
rect 9368 31471 9444 31557
rect 9368 31415 9378 31471
rect 9434 31415 9444 31471
rect 9368 31329 9444 31415
rect 9368 31273 9378 31329
rect 9434 31273 9444 31329
rect 9368 31187 9444 31273
rect 9368 31131 9378 31187
rect 9434 31131 9444 31187
rect 9368 31045 9444 31131
rect 9368 30989 9378 31045
rect 9434 30989 9444 31045
rect 9368 30903 9444 30989
rect 9368 30847 9378 30903
rect 9434 30847 9444 30903
rect 9368 30761 9444 30847
rect 9368 30705 9378 30761
rect 9434 30705 9444 30761
rect 9368 30695 9444 30705
rect 9784 32323 9860 32333
rect 9784 32267 9794 32323
rect 9850 32267 9860 32323
rect 9784 32181 9860 32267
rect 9784 32125 9794 32181
rect 9850 32125 9860 32181
rect 9784 32039 9860 32125
rect 9784 31983 9794 32039
rect 9850 31983 9860 32039
rect 9784 31897 9860 31983
rect 9784 31841 9794 31897
rect 9850 31841 9860 31897
rect 9784 31755 9860 31841
rect 9784 31699 9794 31755
rect 9850 31699 9860 31755
rect 9784 31613 9860 31699
rect 9784 31557 9794 31613
rect 9850 31557 9860 31613
rect 9784 31471 9860 31557
rect 9784 31415 9794 31471
rect 9850 31415 9860 31471
rect 9784 31329 9860 31415
rect 9784 31273 9794 31329
rect 9850 31273 9860 31329
rect 9784 31187 9860 31273
rect 9784 31131 9794 31187
rect 9850 31131 9860 31187
rect 9784 31045 9860 31131
rect 9784 30989 9794 31045
rect 9850 30989 9860 31045
rect 9784 30903 9860 30989
rect 9784 30847 9794 30903
rect 9850 30847 9860 30903
rect 9784 30761 9860 30847
rect 9784 30705 9794 30761
rect 9850 30705 9860 30761
rect 9784 30695 9860 30705
rect 10272 32323 10348 32333
rect 10272 32267 10282 32323
rect 10338 32267 10348 32323
rect 10272 32181 10348 32267
rect 10272 32125 10282 32181
rect 10338 32125 10348 32181
rect 10272 32039 10348 32125
rect 10272 31983 10282 32039
rect 10338 31983 10348 32039
rect 10272 31897 10348 31983
rect 10272 31841 10282 31897
rect 10338 31841 10348 31897
rect 10272 31755 10348 31841
rect 10272 31699 10282 31755
rect 10338 31699 10348 31755
rect 10272 31613 10348 31699
rect 10272 31557 10282 31613
rect 10338 31557 10348 31613
rect 10272 31471 10348 31557
rect 10272 31415 10282 31471
rect 10338 31415 10348 31471
rect 10272 31329 10348 31415
rect 10272 31273 10282 31329
rect 10338 31273 10348 31329
rect 10272 31187 10348 31273
rect 10272 31131 10282 31187
rect 10338 31131 10348 31187
rect 10272 31045 10348 31131
rect 10272 30989 10282 31045
rect 10338 30989 10348 31045
rect 10272 30903 10348 30989
rect 10272 30847 10282 30903
rect 10338 30847 10348 30903
rect 10272 30761 10348 30847
rect 10272 30705 10282 30761
rect 10338 30705 10348 30761
rect 10272 30695 10348 30705
rect 10760 32272 10836 32282
rect 10760 32216 10770 32272
rect 10826 32216 10836 32272
rect 10760 32130 10836 32216
rect 10760 32074 10770 32130
rect 10826 32074 10836 32130
rect 10760 31988 10836 32074
rect 10760 31932 10770 31988
rect 10826 31932 10836 31988
rect 10760 31846 10836 31932
rect 10760 31790 10770 31846
rect 10826 31790 10836 31846
rect 10760 31704 10836 31790
rect 10760 31648 10770 31704
rect 10826 31648 10836 31704
rect 10760 31562 10836 31648
rect 10760 31506 10770 31562
rect 10826 31506 10836 31562
rect 10760 31420 10836 31506
rect 10760 31364 10770 31420
rect 10826 31364 10836 31420
rect 10760 31278 10836 31364
rect 10760 31222 10770 31278
rect 10826 31222 10836 31278
rect 10760 31136 10836 31222
rect 10760 31080 10770 31136
rect 10826 31080 10836 31136
rect 10760 30994 10836 31080
rect 10760 30938 10770 30994
rect 10826 30938 10836 30994
rect 10760 30852 10836 30938
rect 10760 30796 10770 30852
rect 10826 30796 10836 30852
rect 10760 30710 10836 30796
rect 10760 30654 10770 30710
rect 10826 30654 10836 30710
rect 10760 30644 10836 30654
rect 10998 32251 11074 32337
rect 14400 32496 14410 32552
rect 14466 32496 14552 32552
rect 14608 32496 14694 32552
rect 14750 32496 14760 32552
rect 14400 32410 14760 32496
rect 14400 32354 14410 32410
rect 14466 32354 14552 32410
rect 14608 32354 14694 32410
rect 14750 32354 14760 32410
rect 11724 32323 11800 32333
rect 10998 32195 11008 32251
rect 11064 32195 11074 32251
rect 10998 32109 11074 32195
rect 10998 32053 11008 32109
rect 11064 32053 11074 32109
rect 10998 31967 11074 32053
rect 10998 31911 11008 31967
rect 11064 31911 11074 31967
rect 10998 31825 11074 31911
rect 10998 31769 11008 31825
rect 11064 31769 11074 31825
rect 10998 31683 11074 31769
rect 10998 31627 11008 31683
rect 11064 31627 11074 31683
rect 10998 31541 11074 31627
rect 10998 31485 11008 31541
rect 11064 31485 11074 31541
rect 10998 31399 11074 31485
rect 10998 31343 11008 31399
rect 11064 31343 11074 31399
rect 10998 31257 11074 31343
rect 10998 31201 11008 31257
rect 11064 31201 11074 31257
rect 10998 31115 11074 31201
rect 10998 31059 11008 31115
rect 11064 31059 11074 31115
rect 10998 30973 11074 31059
rect 10998 30917 11008 30973
rect 11064 30917 11074 30973
rect 10998 30831 11074 30917
rect 10998 30775 11008 30831
rect 11064 30775 11074 30831
rect 10998 30689 11074 30775
rect 10998 30633 11008 30689
rect 11064 30633 11074 30689
rect 11236 32272 11312 32282
rect 11236 32216 11246 32272
rect 11302 32216 11312 32272
rect 11236 32130 11312 32216
rect 11236 32074 11246 32130
rect 11302 32074 11312 32130
rect 11236 31988 11312 32074
rect 11236 31932 11246 31988
rect 11302 31932 11312 31988
rect 11236 31846 11312 31932
rect 11236 31790 11246 31846
rect 11302 31790 11312 31846
rect 11236 31704 11312 31790
rect 11236 31648 11246 31704
rect 11302 31648 11312 31704
rect 11236 31562 11312 31648
rect 11236 31506 11246 31562
rect 11302 31506 11312 31562
rect 11236 31420 11312 31506
rect 11236 31364 11246 31420
rect 11302 31364 11312 31420
rect 11236 31278 11312 31364
rect 11236 31222 11246 31278
rect 11302 31222 11312 31278
rect 11236 31136 11312 31222
rect 11236 31080 11246 31136
rect 11302 31080 11312 31136
rect 11236 30994 11312 31080
rect 11236 30938 11246 30994
rect 11302 30938 11312 30994
rect 11236 30852 11312 30938
rect 11236 30796 11246 30852
rect 11302 30796 11312 30852
rect 11236 30710 11312 30796
rect 11236 30654 11246 30710
rect 11302 30654 11312 30710
rect 11724 32267 11734 32323
rect 11790 32267 11800 32323
rect 11724 32181 11800 32267
rect 11724 32125 11734 32181
rect 11790 32125 11800 32181
rect 11724 32039 11800 32125
rect 11724 31983 11734 32039
rect 11790 31983 11800 32039
rect 11724 31897 11800 31983
rect 11724 31841 11734 31897
rect 11790 31841 11800 31897
rect 11724 31755 11800 31841
rect 11724 31699 11734 31755
rect 11790 31699 11800 31755
rect 11724 31613 11800 31699
rect 11724 31557 11734 31613
rect 11790 31557 11800 31613
rect 11724 31471 11800 31557
rect 11724 31415 11734 31471
rect 11790 31415 11800 31471
rect 11724 31329 11800 31415
rect 11724 31273 11734 31329
rect 11790 31273 11800 31329
rect 11724 31187 11800 31273
rect 11724 31131 11734 31187
rect 11790 31131 11800 31187
rect 11724 31045 11800 31131
rect 11724 30989 11734 31045
rect 11790 30989 11800 31045
rect 11724 30903 11800 30989
rect 11724 30847 11734 30903
rect 11790 30847 11800 30903
rect 11724 30761 11800 30847
rect 11724 30705 11734 30761
rect 11790 30705 11800 30761
rect 11724 30695 11800 30705
rect 12212 32322 12288 32332
rect 12212 32266 12222 32322
rect 12278 32266 12288 32322
rect 12212 32180 12288 32266
rect 12212 32124 12222 32180
rect 12278 32124 12288 32180
rect 12212 32038 12288 32124
rect 12212 31982 12222 32038
rect 12278 31982 12288 32038
rect 12212 31896 12288 31982
rect 12212 31840 12222 31896
rect 12278 31840 12288 31896
rect 12212 31754 12288 31840
rect 12212 31698 12222 31754
rect 12278 31698 12288 31754
rect 12212 31612 12288 31698
rect 12212 31556 12222 31612
rect 12278 31556 12288 31612
rect 12212 31470 12288 31556
rect 12212 31414 12222 31470
rect 12278 31414 12288 31470
rect 12212 31328 12288 31414
rect 12212 31272 12222 31328
rect 12278 31272 12288 31328
rect 12212 31186 12288 31272
rect 12212 31130 12222 31186
rect 12278 31130 12288 31186
rect 12212 31044 12288 31130
rect 12212 30988 12222 31044
rect 12278 30988 12288 31044
rect 12212 30902 12288 30988
rect 12212 30846 12222 30902
rect 12278 30846 12288 30902
rect 12212 30760 12288 30846
rect 12212 30704 12222 30760
rect 12278 30704 12288 30760
rect 11236 30644 11312 30654
rect 10998 30623 11074 30633
rect 7976 30562 7986 30618
rect 8042 30562 8052 30618
rect 7976 30476 8052 30562
rect 7976 30420 7986 30476
rect 8042 30420 8052 30476
rect 7976 30334 8052 30420
rect 7976 30278 7986 30334
rect 8042 30278 8052 30334
rect 7976 30192 8052 30278
rect 7976 30136 7986 30192
rect 8042 30136 8052 30192
rect 7976 30126 8052 30136
rect 12212 30618 12288 30704
rect 12212 30562 12222 30618
rect 12278 30562 12288 30618
rect 12212 30476 12288 30562
rect 12212 30420 12222 30476
rect 12278 30420 12288 30476
rect 12212 30334 12288 30420
rect 12212 30278 12222 30334
rect 12278 30278 12288 30334
rect 12212 30192 12288 30278
rect 12212 30136 12222 30192
rect 12278 30136 12288 30192
rect 12212 30126 12288 30136
rect 12628 32322 12704 32332
rect 12628 32266 12638 32322
rect 12694 32266 12704 32322
rect 12628 32180 12704 32266
rect 12628 32124 12638 32180
rect 12694 32124 12704 32180
rect 12628 32038 12704 32124
rect 12628 31982 12638 32038
rect 12694 31982 12704 32038
rect 12628 31896 12704 31982
rect 12628 31840 12638 31896
rect 12694 31840 12704 31896
rect 12628 31754 12704 31840
rect 12628 31698 12638 31754
rect 12694 31698 12704 31754
rect 12628 31612 12704 31698
rect 12628 31556 12638 31612
rect 12694 31556 12704 31612
rect 12628 31470 12704 31556
rect 12628 31414 12638 31470
rect 12694 31414 12704 31470
rect 12628 31328 12704 31414
rect 12628 31272 12638 31328
rect 12694 31272 12704 31328
rect 12628 31186 12704 31272
rect 12628 31130 12638 31186
rect 12694 31130 12704 31186
rect 12628 31044 12704 31130
rect 12628 30988 12638 31044
rect 12694 30988 12704 31044
rect 12628 30902 12704 30988
rect 12628 30846 12638 30902
rect 12694 30846 12704 30902
rect 12628 30760 12704 30846
rect 12628 30704 12638 30760
rect 12694 30704 12704 30760
rect 12628 30618 12704 30704
rect 12628 30562 12638 30618
rect 12694 30562 12704 30618
rect 12628 30476 12704 30562
rect 12628 30420 12638 30476
rect 12694 30420 12704 30476
rect 12628 30334 12704 30420
rect 12628 30278 12638 30334
rect 12694 30278 12704 30334
rect 12628 30192 12704 30278
rect 12628 30136 12638 30192
rect 12694 30136 12704 30192
rect 12628 30126 12704 30136
rect 14020 32322 14096 32332
rect 14020 32266 14030 32322
rect 14086 32266 14096 32322
rect 14020 32180 14096 32266
rect 14020 32124 14030 32180
rect 14086 32124 14096 32180
rect 14020 32038 14096 32124
rect 14020 31982 14030 32038
rect 14086 31982 14096 32038
rect 14020 31896 14096 31982
rect 14020 31840 14030 31896
rect 14086 31840 14096 31896
rect 14020 31754 14096 31840
rect 14020 31698 14030 31754
rect 14086 31698 14096 31754
rect 14020 31612 14096 31698
rect 14020 31556 14030 31612
rect 14086 31556 14096 31612
rect 14020 31470 14096 31556
rect 14020 31414 14030 31470
rect 14086 31414 14096 31470
rect 14020 31328 14096 31414
rect 14020 31272 14030 31328
rect 14086 31272 14096 31328
rect 14020 31186 14096 31272
rect 14020 31130 14030 31186
rect 14086 31130 14096 31186
rect 14020 31044 14096 31130
rect 14020 30988 14030 31044
rect 14086 30988 14096 31044
rect 14020 30902 14096 30988
rect 14020 30846 14030 30902
rect 14086 30846 14096 30902
rect 14020 30760 14096 30846
rect 14020 30704 14030 30760
rect 14086 30704 14096 30760
rect 14020 30618 14096 30704
rect 14020 30562 14030 30618
rect 14086 30562 14096 30618
rect 14020 30476 14096 30562
rect 14020 30420 14030 30476
rect 14086 30420 14096 30476
rect 14020 30334 14096 30420
rect 14020 30278 14030 30334
rect 14086 30278 14096 30334
rect 14020 30192 14096 30278
rect 14020 30136 14030 30192
rect 14086 30136 14096 30192
rect 14020 30126 14096 30136
rect 14400 32268 14760 32354
rect 14400 32212 14410 32268
rect 14466 32212 14552 32268
rect 14608 32212 14694 32268
rect 14750 32212 14760 32268
rect 14400 32126 14760 32212
rect 14400 32070 14410 32126
rect 14466 32070 14552 32126
rect 14608 32070 14694 32126
rect 14750 32070 14760 32126
rect 14400 31984 14760 32070
rect 14400 31928 14410 31984
rect 14466 31928 14552 31984
rect 14608 31928 14694 31984
rect 14750 31928 14760 31984
rect 14400 31842 14760 31928
rect 14400 31786 14410 31842
rect 14466 31786 14552 31842
rect 14608 31786 14694 31842
rect 14750 31786 14760 31842
rect 14400 31700 14760 31786
rect 14400 31644 14410 31700
rect 14466 31644 14552 31700
rect 14608 31644 14694 31700
rect 14750 31644 14760 31700
rect 14400 31558 14760 31644
rect 14400 31502 14410 31558
rect 14466 31502 14552 31558
rect 14608 31502 14694 31558
rect 14750 31502 14760 31558
rect 14400 31416 14760 31502
rect 14400 31360 14410 31416
rect 14466 31360 14552 31416
rect 14608 31360 14694 31416
rect 14750 31360 14760 31416
rect 14400 31274 14760 31360
rect 14400 31218 14410 31274
rect 14466 31218 14552 31274
rect 14608 31218 14694 31274
rect 14750 31218 14760 31274
rect 14400 31132 14760 31218
rect 14400 31076 14410 31132
rect 14466 31076 14552 31132
rect 14608 31076 14694 31132
rect 14750 31076 14760 31132
rect 14400 30990 14760 31076
rect 14400 30934 14410 30990
rect 14466 30934 14552 30990
rect 14608 30934 14694 30990
rect 14750 30934 14760 30990
rect 14400 30848 14760 30934
rect 14400 30792 14410 30848
rect 14466 30792 14552 30848
rect 14608 30792 14694 30848
rect 14750 30792 14760 30848
rect 14400 30706 14760 30792
rect 14400 30650 14410 30706
rect 14466 30650 14552 30706
rect 14608 30650 14694 30706
rect 14750 30650 14760 30706
rect 14400 30564 14760 30650
rect 14400 30508 14410 30564
rect 14466 30508 14552 30564
rect 14608 30508 14694 30564
rect 14750 30508 14760 30564
rect 14400 30422 14760 30508
rect 14400 30366 14410 30422
rect 14466 30366 14552 30422
rect 14608 30366 14694 30422
rect 14750 30366 14760 30422
rect 14400 30280 14760 30366
rect 14400 30224 14410 30280
rect 14466 30224 14552 30280
rect 14608 30224 14694 30280
rect 14750 30224 14760 30280
rect 14400 30138 14760 30224
rect 486 30072 562 30082
rect 14400 30082 14410 30138
rect 14466 30082 14552 30138
rect 14608 30082 14694 30138
rect 14750 30082 14760 30138
rect 14400 30072 14760 30082
rect 14400 29797 14760 29807
rect 1985 29739 3339 29749
rect 1985 29683 1995 29739
rect 2051 29683 2137 29739
rect 2193 29683 2279 29739
rect 2335 29683 2421 29739
rect 2477 29683 2563 29739
rect 2619 29683 2705 29739
rect 2761 29683 2847 29739
rect 2903 29683 2989 29739
rect 3045 29683 3131 29739
rect 3187 29683 3273 29739
rect 3329 29683 3339 29739
rect 1985 29673 3339 29683
rect 11922 29739 13276 29749
rect 11922 29683 11932 29739
rect 11988 29683 12074 29739
rect 12130 29683 12216 29739
rect 12272 29683 12358 29739
rect 12414 29683 12500 29739
rect 12556 29683 12642 29739
rect 12698 29683 12784 29739
rect 12840 29683 12926 29739
rect 12982 29683 13068 29739
rect 13124 29683 13210 29739
rect 13266 29683 13276 29739
rect 11922 29673 13276 29683
rect 14400 29741 14410 29797
rect 14466 29741 14552 29797
rect 14608 29741 14694 29797
rect 14750 29741 14760 29797
rect 14400 29655 14760 29741
rect 14400 29599 14410 29655
rect 14466 29599 14552 29655
rect 14608 29599 14694 29655
rect 14750 29599 14760 29655
rect 14400 29513 14760 29599
rect 14400 29457 14410 29513
rect 14466 29457 14552 29513
rect 14608 29457 14694 29513
rect 14750 29457 14760 29513
rect 14400 29371 14760 29457
rect 14400 29315 14410 29371
rect 14466 29315 14552 29371
rect 14608 29315 14694 29371
rect 14750 29315 14760 29371
rect 14400 29229 14760 29315
rect 14400 29173 14410 29229
rect 14466 29173 14552 29229
rect 14608 29173 14694 29229
rect 14750 29173 14760 29229
rect 14400 29087 14760 29173
rect 14400 29031 14410 29087
rect 14466 29031 14552 29087
rect 14608 29031 14694 29087
rect 14750 29031 14760 29087
rect 14400 28945 14760 29031
rect 14400 28889 14410 28945
rect 14466 28889 14552 28945
rect 14608 28889 14694 28945
rect 14750 28889 14760 28945
rect 14400 28803 14760 28889
rect 14400 28747 14410 28803
rect 14466 28747 14552 28803
rect 14608 28747 14694 28803
rect 14750 28747 14760 28803
rect 14400 28661 14760 28747
rect 14400 28605 14410 28661
rect 14466 28605 14552 28661
rect 14608 28605 14694 28661
rect 14750 28605 14760 28661
rect 14400 28519 14760 28605
rect 14400 28463 14410 28519
rect 14466 28463 14552 28519
rect 14608 28463 14694 28519
rect 14750 28463 14760 28519
rect 14400 28453 14760 28463
rect 165 28197 383 28207
rect 165 28141 175 28197
rect 231 28141 317 28197
rect 373 28141 383 28197
rect 165 28055 383 28141
rect 165 27999 175 28055
rect 231 27999 317 28055
rect 373 27999 383 28055
rect 165 27913 383 27999
rect 165 27857 175 27913
rect 231 27857 317 27913
rect 373 27857 383 27913
rect 165 27771 383 27857
rect 165 27715 175 27771
rect 231 27715 317 27771
rect 373 27715 383 27771
rect 165 27629 383 27715
rect 165 27573 175 27629
rect 231 27573 317 27629
rect 373 27573 383 27629
rect 165 27487 383 27573
rect 165 27431 175 27487
rect 231 27431 317 27487
rect 373 27431 383 27487
rect 165 27345 383 27431
rect 165 27289 175 27345
rect 231 27289 317 27345
rect 373 27289 383 27345
rect 165 27203 383 27289
rect 165 27147 175 27203
rect 231 27147 317 27203
rect 373 27147 383 27203
rect 165 27061 383 27147
rect 165 27005 175 27061
rect 231 27005 317 27061
rect 373 27005 383 27061
rect 165 26919 383 27005
rect 165 26863 175 26919
rect 231 26863 317 26919
rect 373 26863 383 26919
rect 165 26853 383 26863
rect 14400 26578 14760 26588
rect 14400 26522 14410 26578
rect 14466 26522 14552 26578
rect 14608 26522 14694 26578
rect 14750 26522 14760 26578
rect 14400 26436 14760 26522
rect 14400 26380 14410 26436
rect 14466 26380 14552 26436
rect 14608 26380 14694 26436
rect 14750 26380 14760 26436
rect 14400 26294 14760 26380
rect 14400 26238 14410 26294
rect 14466 26238 14552 26294
rect 14608 26238 14694 26294
rect 14750 26238 14760 26294
rect 14400 26152 14760 26238
rect 14400 26096 14410 26152
rect 14466 26096 14552 26152
rect 14608 26096 14694 26152
rect 14750 26096 14760 26152
rect 14400 26010 14760 26096
rect 14400 25954 14410 26010
rect 14466 25954 14552 26010
rect 14608 25954 14694 26010
rect 14750 25954 14760 26010
rect 14400 25868 14760 25954
rect 14400 25812 14410 25868
rect 14466 25812 14552 25868
rect 14608 25812 14694 25868
rect 14750 25812 14760 25868
rect 14400 25726 14760 25812
rect 14400 25670 14410 25726
rect 14466 25670 14552 25726
rect 14608 25670 14694 25726
rect 14750 25670 14760 25726
rect 14400 25584 14760 25670
rect 14400 25528 14410 25584
rect 14466 25528 14552 25584
rect 14608 25528 14694 25584
rect 14750 25528 14760 25584
rect 14400 25442 14760 25528
rect 14400 25386 14410 25442
rect 14466 25386 14552 25442
rect 14608 25386 14694 25442
rect 14750 25386 14760 25442
rect 14400 25300 14760 25386
rect 14400 25244 14410 25300
rect 14466 25244 14552 25300
rect 14608 25244 14694 25300
rect 14750 25244 14760 25300
rect 14400 25158 14760 25244
rect 14400 25102 14410 25158
rect 14466 25102 14552 25158
rect 14608 25102 14694 25158
rect 14750 25102 14760 25158
rect 14400 25016 14760 25102
rect 14400 24960 14410 25016
rect 14466 24960 14552 25016
rect 14608 24960 14694 25016
rect 14750 24960 14760 25016
rect 14400 24874 14760 24960
rect 14400 24818 14410 24874
rect 14466 24818 14552 24874
rect 14608 24818 14694 24874
rect 14750 24818 14760 24874
rect 14400 24732 14760 24818
rect 14400 24676 14410 24732
rect 14466 24676 14552 24732
rect 14608 24676 14694 24732
rect 14750 24676 14760 24732
rect 14400 24590 14760 24676
rect 14400 24534 14410 24590
rect 14466 24534 14552 24590
rect 14608 24534 14694 24590
rect 14750 24534 14760 24590
rect 14400 24448 14760 24534
rect 14400 24392 14410 24448
rect 14466 24392 14552 24448
rect 14608 24392 14694 24448
rect 14750 24392 14760 24448
rect 14400 24306 14760 24392
rect 14400 24250 14410 24306
rect 14466 24250 14552 24306
rect 14608 24250 14694 24306
rect 14750 24250 14760 24306
rect 14400 24164 14760 24250
rect 14400 24108 14410 24164
rect 14466 24108 14552 24164
rect 14608 24108 14694 24164
rect 14750 24108 14760 24164
rect 14400 24022 14760 24108
rect 14400 23966 14410 24022
rect 14466 23966 14552 24022
rect 14608 23966 14694 24022
rect 14750 23966 14760 24022
rect 14400 23880 14760 23966
rect 14400 23824 14410 23880
rect 14466 23824 14552 23880
rect 14608 23824 14694 23880
rect 14750 23824 14760 23880
rect 14400 23738 14760 23824
rect 14400 23682 14410 23738
rect 14466 23682 14552 23738
rect 14608 23682 14694 23738
rect 14750 23682 14760 23738
rect 14400 23672 14760 23682
rect 14400 23378 14760 23388
rect 14400 23322 14410 23378
rect 14466 23322 14552 23378
rect 14608 23322 14694 23378
rect 14750 23322 14760 23378
rect 14400 23236 14760 23322
rect 14400 23180 14410 23236
rect 14466 23180 14552 23236
rect 14608 23180 14694 23236
rect 14750 23180 14760 23236
rect 14400 23094 14760 23180
rect 14400 23038 14410 23094
rect 14466 23038 14552 23094
rect 14608 23038 14694 23094
rect 14750 23038 14760 23094
rect 14400 22952 14760 23038
rect 14400 22896 14410 22952
rect 14466 22896 14552 22952
rect 14608 22896 14694 22952
rect 14750 22896 14760 22952
rect 14400 22810 14760 22896
rect 14400 22754 14410 22810
rect 14466 22754 14552 22810
rect 14608 22754 14694 22810
rect 14750 22754 14760 22810
rect 14400 22668 14760 22754
rect 14400 22612 14410 22668
rect 14466 22612 14552 22668
rect 14608 22612 14694 22668
rect 14750 22612 14760 22668
rect 14400 22526 14760 22612
rect 14400 22470 14410 22526
rect 14466 22470 14552 22526
rect 14608 22470 14694 22526
rect 14750 22470 14760 22526
rect 14400 22384 14760 22470
rect 14400 22328 14410 22384
rect 14466 22328 14552 22384
rect 14608 22328 14694 22384
rect 14750 22328 14760 22384
rect 14400 22242 14760 22328
rect 14400 22186 14410 22242
rect 14466 22186 14552 22242
rect 14608 22186 14694 22242
rect 14750 22186 14760 22242
rect 14400 22100 14760 22186
rect 14400 22044 14410 22100
rect 14466 22044 14552 22100
rect 14608 22044 14694 22100
rect 14750 22044 14760 22100
rect 14400 21958 14760 22044
rect 14400 21902 14410 21958
rect 14466 21902 14552 21958
rect 14608 21902 14694 21958
rect 14750 21902 14760 21958
rect 14400 21816 14760 21902
rect 14400 21760 14410 21816
rect 14466 21760 14552 21816
rect 14608 21760 14694 21816
rect 14750 21760 14760 21816
rect 14400 21674 14760 21760
rect 14400 21618 14410 21674
rect 14466 21618 14552 21674
rect 14608 21618 14694 21674
rect 14750 21618 14760 21674
rect 14400 21532 14760 21618
rect 14400 21476 14410 21532
rect 14466 21476 14552 21532
rect 14608 21476 14694 21532
rect 14750 21476 14760 21532
rect 14400 21390 14760 21476
rect 14400 21334 14410 21390
rect 14466 21334 14552 21390
rect 14608 21334 14694 21390
rect 14750 21334 14760 21390
rect 14400 21248 14760 21334
rect 14400 21192 14410 21248
rect 14466 21192 14552 21248
rect 14608 21192 14694 21248
rect 14750 21192 14760 21248
rect 14400 21106 14760 21192
rect 14400 21050 14410 21106
rect 14466 21050 14552 21106
rect 14608 21050 14694 21106
rect 14750 21050 14760 21106
rect 14400 20964 14760 21050
rect 14400 20908 14410 20964
rect 14466 20908 14552 20964
rect 14608 20908 14694 20964
rect 14750 20908 14760 20964
rect 14400 20822 14760 20908
rect 14400 20766 14410 20822
rect 14466 20766 14552 20822
rect 14608 20766 14694 20822
rect 14750 20766 14760 20822
rect 14400 20680 14760 20766
rect 14400 20624 14410 20680
rect 14466 20624 14552 20680
rect 14608 20624 14694 20680
rect 14750 20624 14760 20680
rect 14400 20538 14760 20624
rect 14400 20482 14410 20538
rect 14466 20482 14552 20538
rect 14608 20482 14694 20538
rect 14750 20482 14760 20538
rect 14400 20472 14760 20482
rect 14400 20178 14760 20188
rect 14400 20122 14410 20178
rect 14466 20122 14552 20178
rect 14608 20122 14694 20178
rect 14750 20122 14760 20178
rect 14400 20036 14760 20122
rect 14400 19980 14410 20036
rect 14466 19980 14552 20036
rect 14608 19980 14694 20036
rect 14750 19980 14760 20036
rect 14400 19894 14760 19980
rect 14400 19838 14410 19894
rect 14466 19838 14552 19894
rect 14608 19838 14694 19894
rect 14750 19838 14760 19894
rect 14400 19752 14760 19838
rect 14400 19696 14410 19752
rect 14466 19696 14552 19752
rect 14608 19696 14694 19752
rect 14750 19696 14760 19752
rect 14400 19610 14760 19696
rect 14400 19554 14410 19610
rect 14466 19554 14552 19610
rect 14608 19554 14694 19610
rect 14750 19554 14760 19610
rect 14400 19468 14760 19554
rect 14400 19412 14410 19468
rect 14466 19412 14552 19468
rect 14608 19412 14694 19468
rect 14750 19412 14760 19468
rect 14400 19326 14760 19412
rect 14400 19270 14410 19326
rect 14466 19270 14552 19326
rect 14608 19270 14694 19326
rect 14750 19270 14760 19326
rect 14400 19184 14760 19270
rect 14400 19128 14410 19184
rect 14466 19128 14552 19184
rect 14608 19128 14694 19184
rect 14750 19128 14760 19184
rect 14400 19042 14760 19128
rect 14400 18986 14410 19042
rect 14466 18986 14552 19042
rect 14608 18986 14694 19042
rect 14750 18986 14760 19042
rect 14400 18900 14760 18986
rect 14400 18844 14410 18900
rect 14466 18844 14552 18900
rect 14608 18844 14694 18900
rect 14750 18844 14760 18900
rect 14400 18758 14760 18844
rect 14400 18702 14410 18758
rect 14466 18702 14552 18758
rect 14608 18702 14694 18758
rect 14750 18702 14760 18758
rect 14400 18616 14760 18702
rect 14400 18560 14410 18616
rect 14466 18560 14552 18616
rect 14608 18560 14694 18616
rect 14750 18560 14760 18616
rect 14400 18474 14760 18560
rect 14400 18418 14410 18474
rect 14466 18418 14552 18474
rect 14608 18418 14694 18474
rect 14750 18418 14760 18474
rect 14400 18332 14760 18418
rect 14400 18276 14410 18332
rect 14466 18276 14552 18332
rect 14608 18276 14694 18332
rect 14750 18276 14760 18332
rect 14400 18190 14760 18276
rect 14400 18134 14410 18190
rect 14466 18134 14552 18190
rect 14608 18134 14694 18190
rect 14750 18134 14760 18190
rect 14400 18048 14760 18134
rect 14400 17992 14410 18048
rect 14466 17992 14552 18048
rect 14608 17992 14694 18048
rect 14750 17992 14760 18048
rect 14400 17906 14760 17992
rect 14400 17850 14410 17906
rect 14466 17850 14552 17906
rect 14608 17850 14694 17906
rect 14750 17850 14760 17906
rect 14400 17764 14760 17850
rect 14400 17708 14410 17764
rect 14466 17708 14552 17764
rect 14608 17708 14694 17764
rect 14750 17708 14760 17764
rect 14400 17622 14760 17708
rect 14400 17566 14410 17622
rect 14466 17566 14552 17622
rect 14608 17566 14694 17622
rect 14750 17566 14760 17622
rect 14400 17480 14760 17566
rect 14400 17424 14410 17480
rect 14466 17424 14552 17480
rect 14608 17424 14694 17480
rect 14750 17424 14760 17480
rect 14400 17338 14760 17424
rect 14400 17282 14410 17338
rect 14466 17282 14552 17338
rect 14608 17282 14694 17338
rect 14750 17282 14760 17338
rect 14400 17272 14760 17282
rect 14400 16978 14760 16988
rect 14400 16922 14410 16978
rect 14466 16922 14552 16978
rect 14608 16922 14694 16978
rect 14750 16922 14760 16978
rect 14400 16836 14760 16922
rect 14400 16780 14410 16836
rect 14466 16780 14552 16836
rect 14608 16780 14694 16836
rect 14750 16780 14760 16836
rect 14400 16694 14760 16780
rect 14400 16638 14410 16694
rect 14466 16638 14552 16694
rect 14608 16638 14694 16694
rect 14750 16638 14760 16694
rect 14400 16552 14760 16638
rect 14400 16496 14410 16552
rect 14466 16496 14552 16552
rect 14608 16496 14694 16552
rect 14750 16496 14760 16552
rect 14400 16410 14760 16496
rect 14400 16354 14410 16410
rect 14466 16354 14552 16410
rect 14608 16354 14694 16410
rect 14750 16354 14760 16410
rect 14400 16268 14760 16354
rect 14400 16212 14410 16268
rect 14466 16212 14552 16268
rect 14608 16212 14694 16268
rect 14750 16212 14760 16268
rect 14400 16126 14760 16212
rect 14400 16070 14410 16126
rect 14466 16070 14552 16126
rect 14608 16070 14694 16126
rect 14750 16070 14760 16126
rect 14400 15984 14760 16070
rect 14400 15928 14410 15984
rect 14466 15928 14552 15984
rect 14608 15928 14694 15984
rect 14750 15928 14760 15984
rect 14400 15842 14760 15928
rect 14400 15786 14410 15842
rect 14466 15786 14552 15842
rect 14608 15786 14694 15842
rect 14750 15786 14760 15842
rect 14400 15700 14760 15786
rect 14400 15644 14410 15700
rect 14466 15644 14552 15700
rect 14608 15644 14694 15700
rect 14750 15644 14760 15700
rect 14400 15558 14760 15644
rect 14400 15502 14410 15558
rect 14466 15502 14552 15558
rect 14608 15502 14694 15558
rect 14750 15502 14760 15558
rect 14400 15416 14760 15502
rect 14400 15360 14410 15416
rect 14466 15360 14552 15416
rect 14608 15360 14694 15416
rect 14750 15360 14760 15416
rect 14400 15274 14760 15360
rect 14400 15218 14410 15274
rect 14466 15218 14552 15274
rect 14608 15218 14694 15274
rect 14750 15218 14760 15274
rect 14400 15132 14760 15218
rect 14400 15076 14410 15132
rect 14466 15076 14552 15132
rect 14608 15076 14694 15132
rect 14750 15076 14760 15132
rect 14400 14990 14760 15076
rect 14400 14934 14410 14990
rect 14466 14934 14552 14990
rect 14608 14934 14694 14990
rect 14750 14934 14760 14990
rect 14400 14848 14760 14934
rect 14400 14792 14410 14848
rect 14466 14792 14552 14848
rect 14608 14792 14694 14848
rect 14750 14792 14760 14848
rect 14400 14706 14760 14792
rect 14400 14650 14410 14706
rect 14466 14650 14552 14706
rect 14608 14650 14694 14706
rect 14750 14650 14760 14706
rect 14400 14564 14760 14650
rect 14400 14508 14410 14564
rect 14466 14508 14552 14564
rect 14608 14508 14694 14564
rect 14750 14508 14760 14564
rect 14400 14422 14760 14508
rect 14400 14366 14410 14422
rect 14466 14366 14552 14422
rect 14608 14366 14694 14422
rect 14750 14366 14760 14422
rect 14400 14280 14760 14366
rect 14400 14224 14410 14280
rect 14466 14224 14552 14280
rect 14608 14224 14694 14280
rect 14750 14224 14760 14280
rect 14400 14138 14760 14224
rect 14400 14082 14410 14138
rect 14466 14082 14552 14138
rect 14608 14082 14694 14138
rect 14750 14082 14760 14138
rect 14400 14072 14760 14082
rect 165 10578 383 10588
rect 165 10522 175 10578
rect 231 10522 317 10578
rect 373 10522 383 10578
rect 165 10436 383 10522
rect 165 10380 175 10436
rect 231 10380 317 10436
rect 373 10380 383 10436
rect 165 10294 383 10380
rect 165 10238 175 10294
rect 231 10238 317 10294
rect 373 10238 383 10294
rect 165 10152 383 10238
rect 165 10096 175 10152
rect 231 10096 317 10152
rect 373 10096 383 10152
rect 165 10010 383 10096
rect 165 9954 175 10010
rect 231 9954 317 10010
rect 373 9954 383 10010
rect 165 9868 383 9954
rect 165 9812 175 9868
rect 231 9812 317 9868
rect 373 9812 383 9868
rect 165 9726 383 9812
rect 165 9670 175 9726
rect 231 9670 317 9726
rect 373 9670 383 9726
rect 165 9584 383 9670
rect 165 9528 175 9584
rect 231 9528 317 9584
rect 373 9528 383 9584
rect 165 9442 383 9528
rect 165 9386 175 9442
rect 231 9386 317 9442
rect 373 9386 383 9442
rect 165 9300 383 9386
rect 165 9244 175 9300
rect 231 9244 317 9300
rect 373 9244 383 9300
rect 165 9158 383 9244
rect 165 9102 175 9158
rect 231 9102 317 9158
rect 373 9102 383 9158
rect 165 9016 383 9102
rect 165 8960 175 9016
rect 231 8960 317 9016
rect 373 8960 383 9016
rect 165 8874 383 8960
rect 165 8818 175 8874
rect 231 8818 317 8874
rect 373 8818 383 8874
rect 165 8732 383 8818
rect 165 8676 175 8732
rect 231 8676 317 8732
rect 373 8676 383 8732
rect 165 8590 383 8676
rect 165 8534 175 8590
rect 231 8534 317 8590
rect 373 8534 383 8590
rect 165 8448 383 8534
rect 165 8392 175 8448
rect 231 8392 317 8448
rect 373 8392 383 8448
rect 165 8306 383 8392
rect 165 8250 175 8306
rect 231 8250 317 8306
rect 373 8250 383 8306
rect 165 8164 383 8250
rect 165 8108 175 8164
rect 231 8108 317 8164
rect 373 8108 383 8164
rect 165 8022 383 8108
rect 165 7966 175 8022
rect 231 7966 317 8022
rect 373 7966 383 8022
rect 165 7880 383 7966
rect 165 7824 175 7880
rect 231 7824 317 7880
rect 373 7824 383 7880
rect 165 7738 383 7824
rect 165 7682 175 7738
rect 231 7682 317 7738
rect 373 7682 383 7738
rect 165 7672 383 7682
rect 165 7378 383 7388
rect 165 7322 175 7378
rect 231 7322 317 7378
rect 373 7322 383 7378
rect 165 7236 383 7322
rect 165 7180 175 7236
rect 231 7180 317 7236
rect 373 7180 383 7236
rect 165 7094 383 7180
rect 165 7038 175 7094
rect 231 7038 317 7094
rect 373 7038 383 7094
rect 165 6952 383 7038
rect 165 6896 175 6952
rect 231 6896 317 6952
rect 373 6896 383 6952
rect 165 6810 383 6896
rect 165 6754 175 6810
rect 231 6754 317 6810
rect 373 6754 383 6810
rect 165 6668 383 6754
rect 165 6612 175 6668
rect 231 6612 317 6668
rect 373 6612 383 6668
rect 165 6526 383 6612
rect 165 6470 175 6526
rect 231 6470 317 6526
rect 373 6470 383 6526
rect 165 6384 383 6470
rect 165 6328 175 6384
rect 231 6328 317 6384
rect 373 6328 383 6384
rect 165 6242 383 6328
rect 165 6186 175 6242
rect 231 6186 317 6242
rect 373 6186 383 6242
rect 165 6100 383 6186
rect 165 6044 175 6100
rect 231 6044 317 6100
rect 373 6044 383 6100
rect 165 5958 383 6044
rect 165 5902 175 5958
rect 231 5902 317 5958
rect 373 5902 383 5958
rect 165 5816 383 5902
rect 165 5760 175 5816
rect 231 5760 317 5816
rect 373 5760 383 5816
rect 165 5674 383 5760
rect 165 5618 175 5674
rect 231 5618 317 5674
rect 373 5618 383 5674
rect 165 5532 383 5618
rect 165 5476 175 5532
rect 231 5476 317 5532
rect 373 5476 383 5532
rect 165 5390 383 5476
rect 165 5334 175 5390
rect 231 5334 317 5390
rect 373 5334 383 5390
rect 165 5248 383 5334
rect 165 5192 175 5248
rect 231 5192 317 5248
rect 373 5192 383 5248
rect 165 5106 383 5192
rect 165 5050 175 5106
rect 231 5050 317 5106
rect 373 5050 383 5106
rect 165 4964 383 5050
rect 165 4908 175 4964
rect 231 4908 317 4964
rect 373 4908 383 4964
rect 165 4822 383 4908
rect 165 4766 175 4822
rect 231 4766 317 4822
rect 373 4766 383 4822
rect 165 4680 383 4766
rect 165 4624 175 4680
rect 231 4624 317 4680
rect 373 4624 383 4680
rect 165 4538 383 4624
rect 165 4482 175 4538
rect 231 4482 317 4538
rect 373 4482 383 4538
rect 165 4472 383 4482
rect 165 4178 383 4188
rect 165 4122 175 4178
rect 231 4122 317 4178
rect 373 4122 383 4178
rect 165 4036 383 4122
rect 165 3980 175 4036
rect 231 3980 317 4036
rect 373 3980 383 4036
rect 165 3894 383 3980
rect 165 3838 175 3894
rect 231 3838 317 3894
rect 373 3838 383 3894
rect 165 3752 383 3838
rect 165 3696 175 3752
rect 231 3696 317 3752
rect 373 3696 383 3752
rect 165 3610 383 3696
rect 165 3554 175 3610
rect 231 3554 317 3610
rect 373 3554 383 3610
rect 165 3468 383 3554
rect 165 3412 175 3468
rect 231 3412 317 3468
rect 373 3412 383 3468
rect 165 3326 383 3412
rect 165 3270 175 3326
rect 231 3270 317 3326
rect 373 3270 383 3326
rect 165 3184 383 3270
rect 165 3128 175 3184
rect 231 3128 317 3184
rect 373 3128 383 3184
rect 165 3042 383 3128
rect 165 2986 175 3042
rect 231 2986 317 3042
rect 373 2986 383 3042
rect 165 2900 383 2986
rect 165 2844 175 2900
rect 231 2844 317 2900
rect 373 2844 383 2900
rect 165 2758 383 2844
rect 165 2702 175 2758
rect 231 2702 317 2758
rect 373 2702 383 2758
rect 165 2616 383 2702
rect 165 2560 175 2616
rect 231 2560 317 2616
rect 373 2560 383 2616
rect 165 2474 383 2560
rect 165 2418 175 2474
rect 231 2418 317 2474
rect 373 2418 383 2474
rect 165 2332 383 2418
rect 165 2276 175 2332
rect 231 2276 317 2332
rect 373 2276 383 2332
rect 165 2190 383 2276
rect 165 2134 175 2190
rect 231 2134 317 2190
rect 373 2134 383 2190
rect 165 2048 383 2134
rect 165 1992 175 2048
rect 231 1992 317 2048
rect 373 1992 383 2048
rect 165 1906 383 1992
rect 165 1850 175 1906
rect 231 1850 317 1906
rect 373 1850 383 1906
rect 165 1764 383 1850
rect 165 1708 175 1764
rect 231 1708 317 1764
rect 373 1708 383 1764
rect 165 1622 383 1708
rect 165 1566 175 1622
rect 231 1566 317 1622
rect 373 1566 383 1622
rect 165 1480 383 1566
rect 165 1424 175 1480
rect 231 1424 317 1480
rect 373 1424 383 1480
rect 165 1338 383 1424
rect 165 1282 175 1338
rect 231 1282 317 1338
rect 373 1282 383 1338
rect 165 1272 383 1282
use comp018green_esd_cdm  comp018green_esd_cdm_0
timestamp 1750858719
transform 1 0 4583 0 -1 49089
box -205 -83 5981 8547
use comp018green_inpath_cms_smt  comp018green_inpath_cms_smt_0
timestamp 1750858719
transform 1 0 848 0 -1 55482
box -144 -83 13504 14940
use comp018green_out_paddrv_24T  comp018green_out_paddrv_24T_0
timestamp 1750858719
transform 1 0 794 0 1 1095
box -462 -1095 13938 27676
use comp018green_out_predrv  comp018green_out_predrv_0
timestamp 1750858719
transform 1 0 479 0 -1 35599
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_1
timestamp 1750858719
transform -1 0 14585 0 -1 35599
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_2
timestamp 1750858719
transform 1 0 7487 0 -1 35599
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_3
timestamp 1750858719
transform -1 0 7577 0 -1 35599
box -83 -83 3677 6020
use comp018green_out_sigbuf_a  comp018green_out_sigbuf_a_0
timestamp 1750858719
transform -1 0 11282 0 1 37131
box -83 -83 2701 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_0
timestamp 1750858719
transform 1 0 798 0 1 37131
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_1
timestamp 1750858719
transform -1 0 6132 0 1 37131
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_2
timestamp 1750858719
transform 1 0 6042 0 1 37131
box -83 -803 2795 2911
use comp018green_sigbuf_1  comp018green_sigbuf_1_0
timestamp 1750858719
transform 1 0 11192 0 1 37131
box -83 -83 2889 2911
use M1_NWELL_CDNS_40661956134321  M1_NWELL_CDNS_40661956134321_0
timestamp 1750858719
transform 1 0 2049 0 1 55282
box 0 0 1 1
use M1_NWELL_CDNS_40661956134321  M1_NWELL_CDNS_40661956134321_1
timestamp 1750858719
transform 1 0 1083 0 1 55282
box 0 0 1 1
use M1_NWELL_CDNS_40661956134322  M1_NWELL_CDNS_40661956134322_0
timestamp 1750858719
transform 1 0 1566 0 1 54765
box 0 0 1 1
use M1_NWELL_CDNS_40661956134322  M1_NWELL_CDNS_40661956134322_1
timestamp 1750858719
transform 1 0 1566 0 1 55799
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134271  M1_PACTIVE_CDNS_40661956134271_0
timestamp 1750858719
transform 1 0 14615 0 1 41962
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134271  M1_PACTIVE_CDNS_40661956134271_1
timestamp 1750858719
transform 1 0 12098 0 1 41962
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134272  M1_PACTIVE_CDNS_40661956134272_0
timestamp 1750858719
transform 1 0 13333 0 1 40740
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134272  M1_PACTIVE_CDNS_40661956134272_1
timestamp 1750858719
transform 1 0 13333 0 1 43184
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134273  M1_PACTIVE_CDNS_40661956134273_0
timestamp 1750858719
transform 1 0 2376 0 1 56269
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134273  M1_PACTIVE_CDNS_40661956134273_1
timestamp 1750858719
transform 1 0 14690 0 1 56269
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134274  M1_PACTIVE_CDNS_40661956134274_0
timestamp 1750858719
transform 0 -1 8533 1 0 55729
box 0 0 1 1
use M1_PACTIVE_CDNS_40661956134274  M1_PACTIVE_CDNS_40661956134274_1
timestamp 1750858719
transform 0 -1 8533 1 0 56809
box 0 0 1 1
use M1_PSUB_CDNS_40661956134319  M1_PSUB_CDNS_40661956134319_0
timestamp 1750858719
transform 1 0 11300 0 1 42779
box 0 0 1 1
use M1_PSUB_CDNS_40661956134324  M1_PSUB_CDNS_40661956134324_0
timestamp 1750858719
transform -1 0 14496 0 1 4964
box 0 0 1 1
use M1_PSUB_CDNS_40661956134324  M1_PSUB_CDNS_40661956134324_1
timestamp 1750858719
transform 1 0 550 0 1 4964
box 0 0 1 1
use M2_M1_CDNS_4066195613432  M2_M1_CDNS_4066195613432_0
timestamp 1750858719
transform 1 0 4140 0 1 48332
box 0 0 1 1
use M2_M1_CDNS_40661956134232  M2_M1_CDNS_40661956134232_0
timestamp 1750858719
transform 1 0 6684 0 1 52283
box 0 0 1 1
use M2_M1_CDNS_40661956134234  M2_M1_CDNS_40661956134234_0
timestamp 1750858719
transform 1 0 10941 0 1 37172
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_0
timestamp 1750858719
transform 1 0 2760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_1
timestamp 1750858719
transform 1 0 6760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_2
timestamp 1750858719
transform 1 0 5760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_3
timestamp 1750858719
transform 1 0 5260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_4
timestamp 1750858719
transform 1 0 4260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_5
timestamp 1750858719
transform 1 0 7260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_6
timestamp 1750858719
transform 1 0 3760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_7
timestamp 1750858719
transform 1 0 9760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_8
timestamp 1750858719
transform 1 0 8760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_9
timestamp 1750858719
transform 1 0 10260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_10
timestamp 1750858719
transform 1 0 8260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_11
timestamp 1750858719
transform 1 0 14470 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_12
timestamp 1750858719
transform 1 0 13260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_13
timestamp 1750858719
transform 1 0 12760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_14
timestamp 1750858719
transform 1 0 11760 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_15
timestamp 1750858719
transform 1 0 11260 0 1 56267
box 0 0 1 1
use M2_M1_CDNS_40661956134236  M2_M1_CDNS_40661956134236_0
timestamp 1750858719
transform 1 0 524 0 1 31583
box 0 0 1 1
use M2_M1_CDNS_40661956134236  M2_M1_CDNS_40661956134236_1
timestamp 1750858719
transform 1 0 14540 0 1 31583
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_0
timestamp 1750858719
transform -1 0 5900 0 1 36230
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_1
timestamp 1750858719
transform -1 0 4580 0 1 35686
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_2
timestamp 1750858719
transform -1 0 6656 0 1 35822
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_3
timestamp 1750858719
transform 1 0 5656 0 1 40202
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_4
timestamp 1750858719
transform -1 0 5484 0 1 35958
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_5
timestamp 1750858719
transform -1 0 7143 0 1 40338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_6
timestamp 1750858719
transform -1 0 4927 0 1 40338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_7
timestamp 1750858719
transform -1 0 4551 0 1 36230
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_8
timestamp 1750858719
transform 1 0 6766 0 1 29241
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_9
timestamp 1750858719
transform 1 0 6522 0 1 29421
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_10
timestamp 1750858719
transform -1 0 6144 0 1 36094
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_11
timestamp 1750858719
transform 1 0 1457 0 1 29421
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_12
timestamp 1750858719
transform 1 0 1686 0 1 40202
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_13
timestamp 1750858719
transform 1 0 2003 0 1 40338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_14
timestamp 1750858719
transform 1 0 3181 0 1 36094
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_15
timestamp 1750858719
transform 1 0 1912 0 1 36094
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_16
timestamp 1750858719
transform 1 0 2572 0 1 35958
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_17
timestamp 1750858719
transform 1 0 1400 0 1 35822
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_18
timestamp 1750858719
transform 1 0 3476 0 1 35686
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_19
timestamp 1750858719
transform 1 0 3586 0 1 29034
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_20
timestamp 1750858719
transform 1 0 1637 0 1 29241
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_21
timestamp 1750858719
transform 1 0 3456 0 1 52611
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_22
timestamp 1750858719
transform 1 0 7344 0 1 52283
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_23
timestamp 1750858719
transform -1 0 3749 0 1 36094
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_24
timestamp 1750858719
transform 1 0 3805 0 1 52611
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_25
timestamp 1750858719
transform 1 0 13425 0 1 35686
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_26
timestamp 1750858719
transform 1 0 13898 0 1 40066
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_27
timestamp 1750858719
transform 1 0 13752 0 1 40202
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_28
timestamp 1750858719
transform 1 0 11506 0 1 40202
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_29
timestamp 1750858719
transform 1 0 13152 0 1 36502
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_30
timestamp 1750858719
transform -1 0 11588 0 1 35686
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_31
timestamp 1750858719
transform -1 0 13664 0 1 35822
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_32
timestamp 1750858719
transform -1 0 12596 0 1 35958
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_33
timestamp 1750858719
transform 1 0 13012 0 1 36366
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_34
timestamp 1750858719
transform -1 0 13429 0 1 29241
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_35
timestamp 1750858719
transform -1 0 11480 0 1 29034
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_36
timestamp 1750858719
transform -1 0 13609 0 1 29421
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_37
timestamp 1750858719
transform 0 -1 11558 1 0 38237
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_38
timestamp 1750858719
transform 0 -1 14096 1 0 40390
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_39
timestamp 1750858719
transform 1 0 12074 0 1 40066
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_40
timestamp 1750858719
transform 1 0 9580 0 1 35958
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_41
timestamp 1750858719
transform 1 0 8408 0 1 35822
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_42
timestamp 1750858719
transform 1 0 10484 0 1 35686
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_43
timestamp 1750858719
transform 1 0 10874 0 1 40338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_44
timestamp 1750858719
transform 1 0 8383 0 1 36366
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_45
timestamp 1750858719
transform -1 0 9060 0 1 36230
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_46
timestamp 1750858719
transform 0 -1 8477 1 0 36554
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_47
timestamp 1750858719
transform 0 -1 11175 1 0 40715
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_48
timestamp 1750858719
transform 1 0 10734 0 1 40066
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_49
timestamp 1750858719
transform 1 0 8657 0 1 35550
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_50
timestamp 1750858719
transform 1 0 8786 0 1 29421
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_51
timestamp 1750858719
transform 1 0 8542 0 1 29241
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_52
timestamp 1750858719
transform 1 0 8920 0 1 36094
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_53
timestamp 1750858719
transform 1 0 12515 0 1 43657
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_0
timestamp 1750858719
transform 1 0 84 0 1 37130
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_1
timestamp 1750858719
transform 1 0 3646 0 1 41930
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_2
timestamp 1750858719
transform 1 0 84 0 1 51530
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_3
timestamp 1750858719
transform 1 0 3646 0 1 43530
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_4
timestamp 1750858719
transform 1 0 14980 0 1 37130
box 0 0 1 1
use M2_M1_CDNS_40661956134240  M2_M1_CDNS_40661956134240_5
timestamp 1750858719
transform 1 0 14980 0 1 51530
box 0 0 1 1
use M2_M1_CDNS_40661956134267  M2_M1_CDNS_40661956134267_0
timestamp 1750858719
transform 1 0 13278 0 1 39918
box 0 0 1 1
use M2_M1_CDNS_40661956134269  M2_M1_CDNS_40661956134269_0
timestamp 1750858719
transform 1 0 3275 0 1 45900
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_0
timestamp 1750858719
transform -1 0 4185 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_1
timestamp 1750858719
transform -1 0 5536 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_2
timestamp 1750858719
transform 1 0 5952 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_3
timestamp 1750858719
transform -1 0 5952 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_4
timestamp 1750858719
transform 1 0 4193 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_5
timestamp 1750858719
transform -1 0 4998 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_6
timestamp 1750858719
transform 1 0 6196 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_7
timestamp 1750858719
transform 1 0 2520 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_8
timestamp 1750858719
transform -1 0 3697 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_9
timestamp 1750858719
transform 1 0 1860 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_10
timestamp 1750858719
transform 1 0 2745 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_11
timestamp 1750858719
transform 1 0 3233 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_12
timestamp 1750858719
transform 1 0 2104 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_13
timestamp 1750858719
transform 1 0 1634 0 1 55452
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_14
timestamp 1750858719
transform 1 0 1492 0 1 55452
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_15
timestamp 1750858719
transform 1 0 11543 0 1 41366
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_16
timestamp 1750858719
transform 1 0 13134 0 1 41493
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_17
timestamp 1750858719
transform 1 0 13570 0 1 41493
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_18
timestamp 1750858719
transform 1 0 11558 0 1 40893
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_19
timestamp 1750858719
transform 1 0 13134 0 1 42420
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_20
timestamp 1750858719
transform 1 0 13341 0 1 38229
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_21
timestamp 1750858719
transform 1 0 13477 0 1 37575
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_22
timestamp 1750858719
transform -1 0 12960 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_23
timestamp 1750858719
transform -1 0 13204 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_24
timestamp 1750858719
transform 1 0 13570 0 1 42420
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_25
timestamp 1750858719
transform -1 0 12544 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_26
timestamp 1750858719
transform 1 0 10068 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_27
timestamp 1750858719
transform 1 0 8933 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_28
timestamp 1750858719
transform -1 0 8331 0 1 38240
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_29
timestamp 1750858719
transform 1 0 9112 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_30
timestamp 1750858719
transform 1 0 10682 0 1 38598
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_31
timestamp 1750858719
transform 1 0 9528 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_32
timestamp 1750858719
transform -1 0 8477 0 1 37491
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_33
timestamp 1750858719
transform -1 0 8868 0 1 33987
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_34
timestamp 1750858719
transform -1 0 10873 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_35
timestamp 1750858719
transform 1 0 10926 0 1 38598
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_36
timestamp 1750858719
transform 1 0 9114 0 1 29021
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_37
timestamp 1750858719
transform 1 0 11634 0 1 47530
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_0
timestamp 1750858719
transform 1 0 6316 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_1
timestamp 1750858719
transform 1 0 5952 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_2
timestamp 1750858719
transform 1 0 5464 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_3
timestamp 1750858719
transform 1 0 4976 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_4
timestamp 1750858719
transform 1 0 7292 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_5
timestamp 1750858719
transform 1 0 4796 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_6
timestamp 1750858719
transform 1 0 7472 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_7
timestamp 1750858719
transform 1 0 4200 0 1 53403
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_8
timestamp 1750858719
transform 1 0 6804 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_9
timestamp 1750858719
transform 1 0 10708 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_10
timestamp 1750858719
transform 1 0 11196 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_11
timestamp 1750858719
transform 1 0 11039 0 1 47014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_12
timestamp 1750858719
transform 1 0 10040 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_13
timestamp 1750858719
transform 1 0 10220 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_14
timestamp 1750858719
transform 1 0 8068 0 1 53403
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_15
timestamp 1750858719
transform 1 0 12716 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_16
timestamp 1750858719
transform 1 0 11560 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_17
timestamp 1750858719
transform 1 0 12048 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_18
timestamp 1750858719
transform 1 0 12536 0 1 55014
box 0 0 1 1
use M2_M1_CDNS_40661956134275  M2_M1_CDNS_40661956134275_19
timestamp 1750858719
transform 1 0 13312 0 1 53403
box 0 0 1 1
use M2_M1_CDNS_40661956134277  M2_M1_CDNS_40661956134277_0
timestamp 1750858719
transform 1 0 6134 0 1 54917
box 0 0 1 1
use M2_M1_CDNS_40661956134277  M2_M1_CDNS_40661956134277_1
timestamp 1750858719
transform 1 0 6134 0 1 53455
box 0 0 1 1
use M2_M1_CDNS_40661956134277  M2_M1_CDNS_40661956134277_2
timestamp 1750858719
transform 1 0 11378 0 1 54917
box 0 0 1 1
use M2_M1_CDNS_40661956134277  M2_M1_CDNS_40661956134277_3
timestamp 1750858719
transform 1 0 11378 0 1 53455
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_0
timestamp 1750858719
transform 1 0 7053 0 1 39132
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_1
timestamp 1750858719
transform 1 0 5121 0 1 39132
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_2
timestamp 1750858719
transform 1 0 1809 0 1 39132
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_3
timestamp 1750858719
transform 1 0 5464 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_4
timestamp 1750858719
transform 1 0 5952 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_5
timestamp 1750858719
transform 1 0 6316 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_6
timestamp 1750858719
transform 1 0 6804 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_7
timestamp 1750858719
transform 1 0 7292 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_8
timestamp 1750858719
transform 1 0 7472 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_9
timestamp 1750858719
transform 1 0 4796 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_10
timestamp 1750858719
transform 1 0 4976 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_11
timestamp 1750858719
transform 1 0 10220 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_12
timestamp 1750858719
transform 1 0 10708 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_13
timestamp 1750858719
transform 1 0 11196 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_14
timestamp 1750858719
transform 1 0 10040 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_15
timestamp 1750858719
transform 1 0 12048 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_16
timestamp 1750858719
transform 1 0 12536 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_17
timestamp 1750858719
transform 1 0 12716 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134279  M2_M1_CDNS_40661956134279_18
timestamp 1750858719
transform 1 0 11560 0 1 53346
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_0
timestamp 1750858719
transform 1 0 6087 0 1 38924
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_1
timestamp 1750858719
transform 1 0 6087 0 1 37648
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_2
timestamp 1750858719
transform 1 0 3465 0 1 37648
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_3
timestamp 1750858719
transform 1 0 843 0 1 37648
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_4
timestamp 1750858719
transform 1 0 3508 0 1 53507
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_5
timestamp 1750858719
transform 1 0 3508 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_6
timestamp 1750858719
transform 1 0 3731 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_7
timestamp 1750858719
transform 1 0 4200 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_8
timestamp 1750858719
transform 1 0 8709 0 1 37648
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_9
timestamp 1750858719
transform 1 0 10365 0 1 38924
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_10
timestamp 1750858719
transform 1 0 10820 0 1 48496
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_11
timestamp 1750858719
transform 1 0 8752 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_12
timestamp 1750858719
transform 1 0 9444 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_13
timestamp 1750858719
transform 1 0 8068 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_14
timestamp 1750858719
transform 1 0 8975 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_15
timestamp 1750858719
transform 1 0 8537 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_16
timestamp 1750858719
transform 1 0 8756 0 1 53507
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_17
timestamp 1750858719
transform 1 0 13312 0 1 54965
box 0 0 1 1
use M2_M1_CDNS_40661956134281  M2_M1_CDNS_40661956134281_18
timestamp 1750858719
transform 1 0 11238 0 1 38924
box 0 0 1 1
use M2_M1_CDNS_40661956134282  M2_M1_CDNS_40661956134282_0
timestamp 1750858719
transform 1 0 4794 0 1 48284
box 0 0 1 1
use M2_M1_CDNS_40661956134283  M2_M1_CDNS_40661956134283_0
timestamp 1750858719
transform 1 0 384 0 1 54575
box 0 0 1 1
use M2_M1_CDNS_40661956134283  M2_M1_CDNS_40661956134283_1
timestamp 1750858719
transform 1 0 384 0 1 53675
box 0 0 1 1
use M2_M1_CDNS_40661956134286  M2_M1_CDNS_40661956134286_0
timestamp 1750858719
transform 1 0 384 0 1 39910
box 0 0 1 1
use M2_M1_CDNS_40661956134286  M2_M1_CDNS_40661956134286_1
timestamp 1750858719
transform 1 0 2270 0 1 36230
box 0 0 1 1
use M2_M1_CDNS_40661956134286  M2_M1_CDNS_40661956134286_2
timestamp 1750858719
transform 1 0 904 0 1 52611
box 0 0 1 1
use M2_M1_CDNS_40661956134286  M2_M1_CDNS_40661956134286_3
timestamp 1750858719
transform 1 0 8616 0 1 49873
box 0 0 1 1
use M2_M1_CDNS_40661956134286  M2_M1_CDNS_40661956134286_4
timestamp 1750858719
transform 1 0 7914 0 1 49873
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_0
timestamp 1750858719
transform 1 0 5713 0 1 48898
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_1
timestamp 1750858719
transform 1 0 7914 0 1 48898
box 0 0 1 1
use M2_M1_CDNS_40661956134287  M2_M1_CDNS_40661956134287_2
timestamp 1750858719
transform 1 0 8616 0 1 48898
box 0 0 1 1
use M2_M1_CDNS_40661956134288  M2_M1_CDNS_40661956134288_0
timestamp 1750858719
transform 1 0 4131 0 1 44941
box 0 0 1 1
use M2_M1_CDNS_40661956134289  M2_M1_CDNS_40661956134289_0
timestamp 1750858719
transform 1 0 3646 0 1 46872
box 0 0 1 1
use M2_M1_CDNS_40661956134291  M2_M1_CDNS_40661956134291_0
timestamp 1750858719
transform 1 0 2758 0 1 40674
box 0 0 1 1
use M2_M1_CDNS_40661956134291  M2_M1_CDNS_40661956134291_1
timestamp 1750858719
transform 1 0 8810 0 1 39918
box 0 0 1 1
use M2_M1_CDNS_40661956134293  M2_M1_CDNS_40661956134293_0
timestamp 1750858719
transform 1 0 4028 0 1 31545
box 0 0 1 1
use M2_M1_CDNS_40661956134293  M2_M1_CDNS_40661956134293_1
timestamp 1750858719
transform 1 0 524 0 1 34666
box 0 0 1 1
use M2_M1_CDNS_40661956134293  M2_M1_CDNS_40661956134293_2
timestamp 1750858719
transform 1 0 11036 0 1 31545
box 0 0 1 1
use M2_M1_CDNS_40661956134295  M2_M1_CDNS_40661956134295_0
timestamp 1750858719
transform 1 0 4334 0 1 49873
box 0 0 1 1
use M2_M1_CDNS_40661956134299  M2_M1_CDNS_40661956134299_0
timestamp 1750858719
transform 1 0 4926 0 1 34874
box 0 0 1 1
use M2_M1_CDNS_40661956134299  M2_M1_CDNS_40661956134299_1
timestamp 1750858719
transform 1 0 3130 0 1 34874
box 0 0 1 1
use M2_M1_CDNS_40661956134299  M2_M1_CDNS_40661956134299_2
timestamp 1750858719
transform 1 0 762 0 1 34874
box 0 0 1 1
use M2_M1_CDNS_40661956134299  M2_M1_CDNS_40661956134299_3
timestamp 1750858719
transform 1 0 11934 0 1 34874
box 0 0 1 1
use M2_M1_CDNS_40661956134299  M2_M1_CDNS_40661956134299_4
timestamp 1750858719
transform 1 0 10138 0 1 34874
box 0 0 1 1
use M2_M1_CDNS_40661956134302  M2_M1_CDNS_40661956134302_0
timestamp 1750858719
transform 1 0 4028 0 1 34250
box 0 0 1 1
use M2_M1_CDNS_40661956134302  M2_M1_CDNS_40661956134302_1
timestamp 1750858719
transform 1 0 11036 0 1 34250
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_0
timestamp 1750858719
transform 1 0 7050 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_1
timestamp 1750858719
transform 1 0 2814 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_2
timestamp 1750858719
transform 1 0 2398 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_3
timestamp 1750858719
transform 1 0 1006 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_4
timestamp 1750858719
transform 1 0 12250 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_5
timestamp 1750858719
transform 1 0 12666 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_6
timestamp 1750858719
transform 1 0 14058 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134305  M2_M1_CDNS_40661956134305_7
timestamp 1750858719
transform 1 0 8014 0 1 31202
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_0
timestamp 1750858719
transform 1 0 5658 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_1
timestamp 1750858719
transform 1 0 5242 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_2
timestamp 1750858719
transform 1 0 4754 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_3
timestamp 1750858719
transform 1 0 4266 0 1 31464
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_4
timestamp 1750858719
transform 1 0 3302 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_5
timestamp 1750858719
transform 1 0 3790 0 1 31464
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_6
timestamp 1750858719
transform 1 0 11762 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_7
timestamp 1750858719
transform 1 0 10310 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_8
timestamp 1750858719
transform 1 0 9822 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_9
timestamp 1750858719
transform 1 0 9406 0 1 31514
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_10
timestamp 1750858719
transform 1 0 10798 0 1 31464
box 0 0 1 1
use M2_M1_CDNS_40661956134307  M2_M1_CDNS_40661956134307_11
timestamp 1750858719
transform 1 0 11274 0 1 31464
box 0 0 1 1
use M2_M1_CDNS_40661956134309  M2_M1_CDNS_40661956134309_0
timestamp 1750858719
transform 1 0 2662 0 1 29711
box 0 0 1 1
use M2_M1_CDNS_40661956134309  M2_M1_CDNS_40661956134309_1
timestamp 1750858719
transform 1 0 12599 0 1 29711
box 0 0 1 1
use M2_M1_CDNS_40661956134315  M2_M1_CDNS_40661956134315_0
timestamp 1750858719
transform 1 0 8066 0 1 55898
box 0 0 1 1
use M2_M1_CDNS_40661956134315  M2_M1_CDNS_40661956134315_1
timestamp 1750858719
transform 1 0 8066 0 1 56640
box 0 0 1 1
use M2_M1_CDNS_40661956134318  M2_M1_CDNS_40661956134318_0
timestamp 1750858719
transform 1 0 3459 0 1 39918
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_0
timestamp 1750858719
transform 1 0 4510 0 1 30306
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_1
timestamp 1750858719
transform 1 0 4998 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_2
timestamp 1750858719
transform 1 0 6562 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_3
timestamp 1750858719
transform 1 0 6806 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_4
timestamp 1750858719
transform 1 0 3546 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_5
timestamp 1750858719
transform 1 0 3058 0 1 30306
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_6
timestamp 1750858719
transform 1 0 1738 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_7
timestamp 1750858719
transform 1 0 1494 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_8
timestamp 1750858719
transform -1 0 12006 0 1 30306
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_9
timestamp 1750858719
transform -1 0 13570 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_10
timestamp 1750858719
transform -1 0 13814 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_11
timestamp 1750858719
transform -1 0 11518 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_12
timestamp 1750858719
transform -1 0 10066 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_13
timestamp 1750858719
transform -1 0 10554 0 1 30306
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_14
timestamp 1750858719
transform 1 0 8746 0 1 30126
box 0 0 1 1
use M2_M1_CDNS_40661956134320  M2_M1_CDNS_40661956134320_15
timestamp 1750858719
transform 1 0 8502 0 1 30126
box 0 0 1 1
use M3_M2_CDNS_4066195613427  M3_M2_CDNS_4066195613427_0
timestamp 1750858719
transform 1 0 4140 0 1 48332
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_0
timestamp 1750858719
transform 1 0 4796 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_1
timestamp 1750858719
transform 1 0 4976 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_2
timestamp 1750858719
transform 1 0 4796 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_3
timestamp 1750858719
transform 1 0 7472 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_4
timestamp 1750858719
transform 1 0 7472 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_5
timestamp 1750858719
transform 1 0 5952 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_6
timestamp 1750858719
transform 1 0 5464 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_7
timestamp 1750858719
transform 1 0 6316 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_8
timestamp 1750858719
transform 1 0 7292 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_9
timestamp 1750858719
transform 1 0 6804 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_10
timestamp 1750858719
transform 1 0 6316 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_11
timestamp 1750858719
transform 1 0 5952 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_12
timestamp 1750858719
transform 1 0 5464 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_13
timestamp 1750858719
transform 1 0 4976 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_14
timestamp 1750858719
transform 1 0 6804 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_15
timestamp 1750858719
transform 1 0 7292 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_16
timestamp 1750858719
transform 1 0 11196 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_17
timestamp 1750858719
transform 1 0 10708 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_18
timestamp 1750858719
transform 1 0 11039 0 1 47014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_19
timestamp 1750858719
transform 1 0 10040 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_20
timestamp 1750858719
transform 1 0 10040 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_21
timestamp 1750858719
transform 1 0 10220 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_22
timestamp 1750858719
transform 1 0 11196 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_23
timestamp 1750858719
transform 1 0 10220 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_24
timestamp 1750858719
transform 1 0 10708 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_25
timestamp 1750858719
transform 1 0 12536 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_26
timestamp 1750858719
transform 1 0 12048 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_27
timestamp 1750858719
transform 1 0 11560 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_28
timestamp 1750858719
transform 1 0 12716 0 1 53346
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_29
timestamp 1750858719
transform 1 0 12716 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_30
timestamp 1750858719
transform 1 0 12048 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_31
timestamp 1750858719
transform 1 0 11560 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134276  M3_M2_CDNS_40661956134276_32
timestamp 1750858719
transform 1 0 12536 0 1 55014
box 0 0 1 1
use M3_M2_CDNS_40661956134278  M3_M2_CDNS_40661956134278_0
timestamp 1750858719
transform 1 0 6134 0 1 53360
box 0 0 1 1
use M3_M2_CDNS_40661956134278  M3_M2_CDNS_40661956134278_1
timestamp 1750858719
transform 1 0 6134 0 1 54917
box 0 0 1 1
use M3_M2_CDNS_40661956134278  M3_M2_CDNS_40661956134278_2
timestamp 1750858719
transform 1 0 11378 0 1 53360
box 0 0 1 1
use M3_M2_CDNS_40661956134278  M3_M2_CDNS_40661956134278_3
timestamp 1750858719
transform 1 0 11378 0 1 54917
box 0 0 1 1
use M3_M2_CDNS_40661956134280  M3_M2_CDNS_40661956134280_0
timestamp 1750858719
transform 1 0 11646 0 1 49428
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_0
timestamp 1750858719
transform 1 0 6087 0 1 37130
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_1
timestamp 1750858719
transform 1 0 3646 0 1 41930
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_2
timestamp 1750858719
transform 1 0 84 0 1 37130
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_3
timestamp 1750858719
transform 1 0 1924 0 1 53130
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_4
timestamp 1750858719
transform 1 0 3646 0 1 43530
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_5
timestamp 1750858719
transform 1 0 84 0 1 51530
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_6
timestamp 1750858719
transform 1 0 14980 0 1 37130
box 0 0 1 1
use M3_M2_CDNS_40661956134284  M3_M2_CDNS_40661956134284_7
timestamp 1750858719
transform 1 0 14980 0 1 51530
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_0
timestamp 1750858719
transform 1 0 384 0 1 38730
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_1
timestamp 1750858719
transform 1 0 904 0 1 37130
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_2
timestamp 1750858719
transform 1 0 384 0 1 49930
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_3
timestamp 1750858719
transform 1 0 904 0 1 51530
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_4
timestamp 1750858719
transform 1 0 14580 0 1 40330
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_5
timestamp 1750858719
transform 1 0 14580 0 1 41930
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_6
timestamp 1750858719
transform 1 0 14580 0 1 29130
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_7
timestamp 1750858719
transform 1 0 9349 0 1 53130
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_8
timestamp 1750858719
transform 1 0 14580 0 1 43530
box 0 0 1 1
use M3_M2_CDNS_40661956134285  M3_M2_CDNS_40661956134285_9
timestamp 1750858719
transform 1 0 14580 0 1 54730
box 0 0 1 1
use M3_M2_CDNS_40661956134290  M3_M2_CDNS_40661956134290_0
timestamp 1750858719
transform 1 0 6087 0 1 38889
box 0 0 1 1
use M3_M2_CDNS_40661956134290  M3_M2_CDNS_40661956134290_1
timestamp 1750858719
transform 1 0 3646 0 1 46889
box 0 0 1 1
use M3_M2_CDNS_40661956134290  M3_M2_CDNS_40661956134290_2
timestamp 1750858719
transform 1 0 10365 0 1 38889
box 0 0 1 1
use M3_M2_CDNS_40661956134290  M3_M2_CDNS_40661956134290_3
timestamp 1750858719
transform 1 0 10820 0 1 48489
box 0 0 1 1
use M3_M2_CDNS_40661956134290  M3_M2_CDNS_40661956134290_4
timestamp 1750858719
transform 1 0 11238 0 1 38889
box 0 0 1 1
use M3_M2_CDNS_40661956134292  M3_M2_CDNS_40661956134292_0
timestamp 1750858719
transform 1 0 2797 0 1 40674
box 0 0 1 1
use M3_M2_CDNS_40661956134294  M3_M2_CDNS_40661956134294_0
timestamp 1750858719
transform 1 0 7053 0 1 39108
box 0 0 1 1
use M3_M2_CDNS_40661956134294  M3_M2_CDNS_40661956134294_1
timestamp 1750858719
transform 1 0 5121 0 1 39108
box 0 0 1 1
use M3_M2_CDNS_40661956134294  M3_M2_CDNS_40661956134294_2
timestamp 1750858719
transform 1 0 1809 0 1 39108
box 0 0 1 1
use M3_M2_CDNS_40661956134296  M3_M2_CDNS_40661956134296_0
timestamp 1750858719
transform 1 0 3460 0 1 39918
box 0 0 1 1
use M3_M2_CDNS_40661956134297  M3_M2_CDNS_40661956134297_0
timestamp 1750858719
transform 1 0 8877 0 1 39918
box 0 0 1 1
use M3_M2_CDNS_40661956134298  M3_M2_CDNS_40661956134298_0
timestamp 1750858719
transform 1 0 13283 0 1 39918
box 0 0 1 1
use M3_M2_CDNS_40661956134298  M3_M2_CDNS_40661956134298_1
timestamp 1750858719
transform 1 0 10960 0 1 37172
box 0 0 1 1
use M3_M2_CDNS_40661956134300  M3_M2_CDNS_40661956134300_0
timestamp 1750858719
transform 1 0 4028 0 1 31584
box 0 0 1 1
use M3_M2_CDNS_40661956134300  M3_M2_CDNS_40661956134300_1
timestamp 1750858719
transform 1 0 524 0 1 34666
box 0 0 1 1
use M3_M2_CDNS_40661956134300  M3_M2_CDNS_40661956134300_2
timestamp 1750858719
transform 1 0 11036 0 1 31584
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_0
timestamp 1750858719
transform 1 0 4926 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_1
timestamp 1750858719
transform 1 0 3130 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_2
timestamp 1750858719
transform 1 0 762 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_3
timestamp 1750858719
transform 1 0 11934 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_4
timestamp 1750858719
transform 1 0 8709 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134301  M3_M2_CDNS_40661956134301_5
timestamp 1750858719
transform 1 0 10138 0 1 34874
box 0 0 1 1
use M3_M2_CDNS_40661956134303  M3_M2_CDNS_40661956134303_0
timestamp 1750858719
transform 1 0 4028 0 1 34481
box 0 0 1 1
use M3_M2_CDNS_40661956134303  M3_M2_CDNS_40661956134303_1
timestamp 1750858719
transform 1 0 11036 0 1 34481
box 0 0 1 1
use M3_M2_CDNS_40661956134304  M3_M2_CDNS_40661956134304_0
timestamp 1750858719
transform 1 0 524 0 1 31530
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_0
timestamp 1750858719
transform 1 0 7050 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_1
timestamp 1750858719
transform 1 0 1006 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_2
timestamp 1750858719
transform 1 0 2814 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_3
timestamp 1750858719
transform 1 0 2398 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_4
timestamp 1750858719
transform 1 0 14058 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_5
timestamp 1750858719
transform 1 0 12666 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_6
timestamp 1750858719
transform 1 0 12250 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134306  M3_M2_CDNS_40661956134306_7
timestamp 1750858719
transform 1 0 8014 0 1 31229
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_0
timestamp 1750858719
transform 1 0 4266 0 1 31463
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_1
timestamp 1750858719
transform 1 0 4754 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_2
timestamp 1750858719
transform 1 0 5242 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_3
timestamp 1750858719
transform 1 0 5658 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_4
timestamp 1750858719
transform 1 0 3302 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_5
timestamp 1750858719
transform 1 0 3790 0 1 31463
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_6
timestamp 1750858719
transform 1 0 11762 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_7
timestamp 1750858719
transform 1 0 9406 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_8
timestamp 1750858719
transform 1 0 9822 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_9
timestamp 1750858719
transform 1 0 10310 0 1 31514
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_10
timestamp 1750858719
transform 1 0 10798 0 1 31463
box 0 0 1 1
use M3_M2_CDNS_40661956134308  M3_M2_CDNS_40661956134308_11
timestamp 1750858719
transform 1 0 11274 0 1 31463
box 0 0 1 1
use M3_M2_CDNS_40661956134310  M3_M2_CDNS_40661956134310_0
timestamp 1750858719
transform 1 0 2662 0 1 29711
box 0 0 1 1
use M3_M2_CDNS_40661956134310  M3_M2_CDNS_40661956134310_1
timestamp 1750858719
transform 1 0 12599 0 1 29711
box 0 0 1 1
use M3_M2_CDNS_40661956134311  M3_M2_CDNS_40661956134311_0
timestamp 1750858719
transform 1 0 14580 0 1 18730
box 0 0 1 1
use M3_M2_CDNS_40661956134311  M3_M2_CDNS_40661956134311_1
timestamp 1750858719
transform 1 0 14580 0 1 25130
box 0 0 1 1
use M3_M2_CDNS_40661956134311  M3_M2_CDNS_40661956134311_2
timestamp 1750858719
transform 1 0 14580 0 1 15530
box 0 0 1 1
use M3_M2_CDNS_40661956134311  M3_M2_CDNS_40661956134311_3
timestamp 1750858719
transform 1 0 14580 0 1 21930
box 0 0 1 1
use M3_M2_CDNS_40661956134311  M3_M2_CDNS_40661956134311_4
timestamp 1750858719
transform 1 0 14580 0 1 31530
box 0 0 1 1
use M3_M2_CDNS_40661956134312  M3_M2_CDNS_40661956134312_0
timestamp 1750858719
transform 1 0 274 0 1 9130
box 0 0 1 1
use M3_M2_CDNS_40661956134312  M3_M2_CDNS_40661956134312_1
timestamp 1750858719
transform 1 0 274 0 1 5930
box 0 0 1 1
use M3_M2_CDNS_40661956134312  M3_M2_CDNS_40661956134312_2
timestamp 1750858719
transform 1 0 274 0 1 2730
box 0 0 1 1
use M3_M2_CDNS_40661956134312  M3_M2_CDNS_40661956134312_3
timestamp 1750858719
transform 1 0 274 0 1 34730
box 0 0 1 1
use M3_M2_CDNS_40661956134313  M3_M2_CDNS_40661956134313_0
timestamp 1750858719
transform 1 0 274 0 1 27530
box 0 0 1 1
use M3_M2_CDNS_40661956134313  M3_M2_CDNS_40661956134313_1
timestamp 1750858719
transform 1 0 12515 0 1 37130
box 0 0 1 1
use M3_M2_CDNS_40661956134314  M3_M2_CDNS_40661956134314_0
timestamp 1750858719
transform 1 0 1924 0 1 56269
box 0 0 1 1
use M3_M2_CDNS_40661956134316  M3_M2_CDNS_40661956134316_0
timestamp 1750858719
transform 1 0 8066 0 1 55898
box 0 0 1 1
use M3_M2_CDNS_40661956134316  M3_M2_CDNS_40661956134316_1
timestamp 1750858719
transform 1 0 8066 0 1 56640
box 0 0 1 1
use M3_M2_CDNS_40661956134317  M3_M2_CDNS_40661956134317_0
timestamp 1750858719
transform 1 0 13331 0 1 42010
box 0 0 1 1
use M3_M2_CDNS_40661956134323  M3_M2_CDNS_40661956134323_0
timestamp 1750858719
transform 1 0 4131 0 1 44941
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613422  nmoscap_6p0_CDNS_4066195613422_0
timestamp 1750858719
transform 0 1 13622 1 0 41178
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613422  nmoscap_6p0_CDNS_4066195613422_1
timestamp 1750858719
transform 0 1 12482 1 0 41178
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613422  nmoscap_6p0_CDNS_4066195613422_2
timestamp 1750858719
transform 0 1 12482 1 0 42146
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613422  nmoscap_6p0_CDNS_4066195613422_3
timestamp 1750858719
transform 0 1 13622 1 0 42146
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_0
timestamp 1750858719
transform 0 1 4260 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_1
timestamp 1750858719
transform 0 1 5760 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_2
timestamp 1750858719
transform 0 1 2760 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_3
timestamp 1750858719
transform 0 1 8760 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_4
timestamp 1750858719
transform 0 1 11760 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_5
timestamp 1750858719
transform 0 1 13260 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_6
timestamp 1750858719
transform 0 1 10260 1 0 56119
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195613423  nmoscap_6p0_CDNS_4066195613423_7
timestamp 1750858719
transform 0 1 7260 1 0 56119
box 0 0 1 1
use pn_6p0_CDNS_4066195613428  pn_6p0_CDNS_4066195613428_0
timestamp 1750858719
transform 1 0 11458 0 1 40793
box 0 0 1 1
use pn_6p0_CDNS_4066195613428  pn_6p0_CDNS_4066195613428_1
timestamp 1750858719
transform 1 0 11458 0 1 41257
box 0 0 1 1
use ppolyf_u_CDNS_4066195613424  ppolyf_u_CDNS_4066195613424_0
timestamp 1750858719
transform 0 -1 1786 1 0 55020
box 0 0 1 1
use ppolyf_u_CDNS_4066195613424  ppolyf_u_CDNS_4066195613424_1
timestamp 1750858719
transform 0 -1 1506 1 0 55020
box 0 0 1 1
<< labels >>
rlabel metal2 s 2136 57117 2136 57117 4 PD
port 1 nsew
rlabel metal2 s 2347 57149 2347 57149 4 IE
port 2 nsew
rlabel metal2 s 7532 28147 7532 28147 4 PAD
port 3 nsew
rlabel metal2 s 13804 57127 13804 57127 4 SL
port 4 nsew
rlabel metal2 s 13950 57170 13950 57170 4 A
port 5 nsew
rlabel metal2 s 14096 57121 14096 57121 4 OE
port 6 nsew
rlabel metal2 s 742 57126 742 57126 4 CS
port 7 nsew
rlabel metal2 s 1263 57113 1263 57113 4 PU
port 8 nsew
rlabel metal2 s 14242 57128 14242 57128 4 Y
port 9 nsew
<< properties >>
string GDS_END 2009696
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1973860
string path 368.350 425.750 368.350 271.325 
<< end >>
