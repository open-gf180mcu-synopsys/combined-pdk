VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_ip_sram__sram512x8m8wm1
  CLASS BLOCK ;
  FOREIGN gf180mcu_fd_ip_sram__sram512x8m8wm1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 431.860 BY 484.880 ;
  SYMMETRY X Y R90 ;
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 145.030 0.000 146.150 5.000 ;
    END
  END A[8]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.525 0.000 149.645 5.000 ;
    END
  END A[7]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 268.860 0.000 269.980 5.000 ;
    END
  END A[6]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 272.085 0.000 273.205 5.000 ;
    END
  END A[5]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 275.820 0.000 276.940 5.000 ;
    END
  END A[4]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 281.325 0.000 282.445 5.000 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.295 0.000 155.415 5.000 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.760 0.000 163.880 5.000 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.215 0.000 172.335 5.000 ;
    END
  END A[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.997600 ;
    PORT
      LAYER Metal2 ;
        RECT 251.710 0.000 252.830 5.000 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 44.706600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.680 0.000 140.800 5.000 ;
    END
  END CLK
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 416.860 0.000 417.980 5.000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 365.150 0.000 366.270 5.000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 358.910 0.000 360.030 5.000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 307.235 0.000 308.355 5.000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.975 0.000 120.095 5.000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.270 0.000 68.390 5.000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.030 0.000 62.150 5.000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.320 0.000 10.440 5.000 ;
    END
  END D[0]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 14.466000 ;
    PORT
      LAYER Metal2 ;
        RECT 202.940 0.000 204.060 5.000 ;
    END
  END GWEN
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 409.275 0.000 410.395 5.000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 368.515 0.000 369.635 5.000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 355.545 0.000 356.665 5.000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 314.790 0.000 315.910 5.000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.395 0.000 112.515 5.000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.635 0.000 71.755 5.000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.665 0.000 58.785 5.000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.328000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.900 0.000 18.020 5.000 ;
    END
  END Q[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 3.530 479.880 428.330 480.880 ;
        RECT 3.530 5.000 5.000 479.880 ;
        RECT 426.860 5.000 428.330 479.880 ;
        RECT 3.530 1.410 8.530 5.000 ;
        RECT 423.330 1.410 428.330 5.000 ;
      LAYER Metal3 ;
        RECT 7.005 480.880 12.005 484.880 ;
        RECT 20.685 480.880 25.685 484.880 ;
        RECT 34.005 480.880 39.005 484.880 ;
        RECT 47.685 480.880 52.685 484.880 ;
        RECT 61.005 480.880 66.005 484.880 ;
        RECT 74.685 480.880 79.685 484.880 ;
        RECT 88.005 480.880 93.005 484.880 ;
        RECT 103.265 480.880 108.265 484.880 ;
        RECT 117.415 480.880 122.415 484.880 ;
        RECT 132.860 480.880 137.860 484.880 ;
        RECT 153.550 480.880 158.550 484.880 ;
        RECT 177.075 480.880 182.075 484.880 ;
        RECT 192.925 480.880 197.925 484.880 ;
        RECT 206.150 480.880 211.150 484.880 ;
        RECT 225.345 480.880 230.345 484.880 ;
        RECT 231.565 480.880 236.565 484.880 ;
        RECT 244.505 480.880 249.505 484.880 ;
        RECT 262.845 480.880 267.845 484.880 ;
        RECT 271.310 480.880 276.310 484.880 ;
        RECT 287.735 480.880 292.735 484.880 ;
        RECT 304.885 480.880 309.885 484.880 ;
        RECT 318.565 480.880 323.565 484.880 ;
        RECT 331.885 480.880 336.885 484.880 ;
        RECT 345.565 480.880 350.565 484.880 ;
        RECT 358.885 480.880 363.885 484.880 ;
        RECT 372.565 480.880 377.565 484.880 ;
        RECT 385.885 480.880 390.885 484.880 ;
        RECT 401.145 480.880 406.145 484.880 ;
        RECT 415.295 480.880 420.295 484.880 ;
        RECT 423.330 480.880 428.330 484.880 ;
        RECT 0.000 479.880 431.860 480.880 ;
        RECT 0.000 475.880 5.000 479.880 ;
        RECT 426.860 475.880 431.860 479.880 ;
        RECT 0.000 466.880 8.530 470.380 ;
        RECT 426.860 466.880 431.860 470.380 ;
        RECT 0.000 457.880 5.000 461.380 ;
        RECT 426.860 457.880 431.860 461.380 ;
        RECT 0.000 448.880 5.000 452.380 ;
        RECT 426.860 448.880 431.860 452.380 ;
        RECT 0.000 439.880 5.000 443.380 ;
        RECT 426.860 439.880 431.860 443.380 ;
        RECT 0.000 430.880 5.000 434.380 ;
        RECT 426.860 430.880 431.860 434.380 ;
        RECT 0.000 421.880 5.000 425.380 ;
        RECT 426.860 421.880 431.860 425.380 ;
        RECT 0.000 412.880 5.000 416.380 ;
        RECT 426.860 412.880 431.860 416.380 ;
        RECT 0.000 403.880 5.000 407.380 ;
        RECT 426.860 403.880 431.860 407.380 ;
        RECT 0.000 394.880 5.000 398.380 ;
        RECT 426.860 394.880 431.860 398.380 ;
        RECT 0.000 385.880 5.000 389.380 ;
        RECT 426.860 385.880 431.860 389.380 ;
        RECT 0.000 376.880 5.000 380.380 ;
        RECT 426.860 376.880 431.860 380.380 ;
        RECT 0.000 367.880 5.000 371.380 ;
        RECT 426.860 367.880 431.860 371.380 ;
        RECT 0.000 358.880 5.000 362.380 ;
        RECT 426.860 358.880 431.860 362.380 ;
        RECT 0.000 349.880 5.000 353.380 ;
        RECT 426.860 349.880 431.860 353.380 ;
        RECT 0.000 340.880 5.000 344.380 ;
        RECT 426.860 340.880 431.860 344.380 ;
        RECT 0.000 331.880 5.000 335.380 ;
        RECT 426.860 331.880 431.860 335.380 ;
        RECT 0.000 322.880 5.000 326.380 ;
        RECT 426.860 322.880 431.860 326.380 ;
        RECT 0.000 313.880 5.000 317.380 ;
        RECT 426.860 313.880 431.860 317.380 ;
        RECT 0.000 304.880 5.000 308.380 ;
        RECT 426.860 304.880 431.860 308.380 ;
        RECT 0.000 295.880 5.000 299.380 ;
        RECT 426.860 295.880 431.860 299.380 ;
        RECT 0.000 286.880 5.000 290.380 ;
        RECT 426.860 286.880 431.860 290.380 ;
        RECT 0.000 277.880 5.000 281.380 ;
        RECT 426.860 277.880 431.860 281.380 ;
        RECT 0.000 268.880 5.000 272.380 ;
        RECT 426.860 268.880 431.860 272.380 ;
        RECT 0.000 259.880 5.000 263.380 ;
        RECT 426.860 259.880 431.860 263.380 ;
        RECT 0.000 250.880 5.000 254.380 ;
        RECT 426.860 250.880 431.860 254.380 ;
        RECT 0.000 241.880 5.000 245.380 ;
        RECT 426.860 241.880 431.860 245.380 ;
        RECT 0.000 232.880 5.000 236.380 ;
        RECT 426.860 232.880 431.860 236.380 ;
        RECT 0.000 223.880 5.000 227.380 ;
        RECT 426.860 223.880 431.860 227.380 ;
        RECT 0.000 214.880 5.000 218.380 ;
        RECT 426.860 214.880 431.860 218.380 ;
        RECT 0.000 205.880 5.000 209.380 ;
        RECT 426.860 205.880 431.860 209.380 ;
        RECT 0.000 196.880 5.000 200.380 ;
        RECT 426.860 196.880 431.860 200.380 ;
        RECT 0.000 187.880 5.000 191.380 ;
        RECT 426.860 187.880 431.860 191.380 ;
        RECT 0.000 178.880 5.000 182.380 ;
        RECT 426.860 178.880 431.860 182.380 ;
        RECT 0.000 147.150 5.000 170.625 ;
        RECT 426.860 147.150 431.860 170.625 ;
        RECT 0.000 114.690 5.000 119.690 ;
        RECT 426.860 114.690 431.860 119.690 ;
        RECT 0.000 90.080 5.000 103.695 ;
        RECT 426.860 90.080 431.860 103.695 ;
        RECT 0.000 60.180 5.000 70.890 ;
        RECT 426.860 60.180 431.860 70.890 ;
        RECT 0.000 40.760 5.000 47.575 ;
        RECT 426.860 40.760 431.860 47.575 ;
        RECT 0.000 20.300 5.000 28.145 ;
        RECT 426.860 20.300 431.860 28.145 ;
        RECT 0.000 6.160 5.000 11.160 ;
        RECT 3.530 5.000 5.000 6.160 ;
        RECT 426.860 6.160 431.860 11.160 ;
        RECT 426.860 5.000 428.330 6.160 ;
        RECT 3.530 0.000 8.530 5.000 ;
        RECT 10.195 0.000 15.195 5.000 ;
        RECT 17.210 0.000 22.210 5.000 ;
        RECT 29.210 0.000 34.210 5.000 ;
        RECT 35.210 0.000 40.210 5.000 ;
        RECT 41.210 0.000 46.210 5.000 ;
        RECT 53.210 0.000 58.210 5.000 ;
        RECT 62.215 0.000 67.215 5.000 ;
        RECT 71.210 0.000 76.210 5.000 ;
        RECT 83.210 0.000 88.210 5.000 ;
        RECT 89.210 0.000 94.210 5.000 ;
        RECT 95.210 0.000 100.210 5.000 ;
        RECT 109.550 0.000 114.550 5.000 ;
        RECT 115.550 0.000 120.550 5.000 ;
        RECT 122.050 0.000 127.050 5.000 ;
        RECT 128.550 0.000 133.550 5.000 ;
        RECT 135.050 0.000 140.050 5.000 ;
        RECT 141.550 0.000 146.550 5.000 ;
        RECT 148.050 0.000 153.050 5.000 ;
        RECT 180.155 0.000 185.155 5.000 ;
        RECT 196.140 0.000 201.140 5.000 ;
        RECT 212.165 0.000 217.165 5.000 ;
        RECT 224.165 0.000 229.165 5.000 ;
        RECT 236.165 0.000 241.165 5.000 ;
        RECT 242.830 0.000 247.830 5.000 ;
        RECT 249.380 0.000 254.380 5.000 ;
        RECT 272.290 0.000 277.290 5.000 ;
        RECT 278.790 0.000 283.790 5.000 ;
        RECT 285.290 0.000 290.290 5.000 ;
        RECT 291.790 0.000 296.790 5.000 ;
        RECT 298.290 0.000 303.290 5.000 ;
        RECT 304.790 0.000 309.790 5.000 ;
        RECT 311.475 0.000 316.475 5.000 ;
        RECT 327.090 0.000 332.090 5.000 ;
        RECT 333.090 0.000 338.090 5.000 ;
        RECT 339.090 0.000 344.090 5.000 ;
        RECT 351.090 0.000 356.090 5.000 ;
        RECT 360.085 0.000 365.085 5.000 ;
        RECT 369.090 0.000 374.090 5.000 ;
        RECT 381.090 0.000 386.090 5.000 ;
        RECT 387.090 0.000 392.090 5.000 ;
        RECT 393.090 0.000 398.090 5.000 ;
        RECT 405.090 0.000 410.090 5.000 ;
        RECT 412.095 0.000 417.095 5.000 ;
        RECT 423.330 0.000 428.330 5.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.130 40.770 143.645 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.685 33.720 173.110 38.260 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.475 161.575 10.940 170.630 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.860 157.430 291.755 160.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.860 136.910 291.755 150.525 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.265 161.575 361.915 170.625 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 133.850 116.850 291.740 121.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.565 99.845 278.225 108.125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 90.075 418.815 103.695 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 119.105 60.230 173.805 64.235 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 251.140 60.175 292.105 69.330 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 299.130 60.175 300.130 70.085 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.035 67.305 362.145 70.890 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 415.845 60.175 421.105 64.235 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 415.845 67.305 421.105 70.895 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 40.770 311.390 47.580 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 363.010 40.760 416.170 47.575 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.435 25.875 136.070 28.150 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 119.545 20.830 312.145 23.095 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 289.545 25.875 312.145 28.150 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.410 479.880 430.450 483.470 ;
        RECT 1.410 5.000 5.000 479.880 ;
        RECT 426.860 5.000 430.450 479.880 ;
        RECT 1.410 1.410 430.450 5.000 ;
      LAYER Metal2 ;
        RECT 1.410 481.840 430.450 483.470 ;
        RECT 1.410 471.390 3.030 474.870 ;
        RECT 428.830 471.390 430.450 474.870 ;
        RECT 1.410 462.390 3.030 465.870 ;
        RECT 428.830 462.390 430.450 465.870 ;
        RECT 1.410 453.390 3.030 456.870 ;
        RECT 428.830 453.390 430.450 456.870 ;
        RECT 1.410 444.390 3.030 447.870 ;
        RECT 428.830 444.390 430.450 447.870 ;
        RECT 1.410 435.390 3.030 438.870 ;
        RECT 428.830 435.390 430.450 438.870 ;
        RECT 1.410 426.390 3.030 429.870 ;
        RECT 428.830 426.390 430.450 429.870 ;
        RECT 1.410 417.390 3.030 420.870 ;
        RECT 428.830 417.390 430.450 420.870 ;
        RECT 1.410 408.390 3.030 411.870 ;
        RECT 428.830 408.390 430.450 411.870 ;
        RECT 1.410 399.390 3.030 402.870 ;
        RECT 428.830 399.390 430.450 402.870 ;
        RECT 1.410 390.390 3.030 393.870 ;
        RECT 428.830 390.390 430.450 393.870 ;
        RECT 1.410 381.390 3.030 384.870 ;
        RECT 428.830 381.390 430.450 384.870 ;
        RECT 1.410 372.390 3.030 375.870 ;
        RECT 428.830 372.390 430.450 375.870 ;
        RECT 1.410 363.390 3.030 366.870 ;
        RECT 428.830 363.390 430.450 366.870 ;
        RECT 1.410 354.390 3.030 357.870 ;
        RECT 428.830 354.390 430.450 357.870 ;
        RECT 1.410 345.390 3.030 348.870 ;
        RECT 428.830 345.390 430.450 348.870 ;
        RECT 1.410 336.390 3.030 339.870 ;
        RECT 428.830 336.390 430.450 339.870 ;
        RECT 1.410 327.390 3.030 330.870 ;
        RECT 428.830 327.390 430.450 330.870 ;
        RECT 1.410 318.390 3.030 321.870 ;
        RECT 428.830 318.390 430.450 321.870 ;
        RECT 1.410 309.390 3.030 312.870 ;
        RECT 428.830 309.390 430.450 312.870 ;
        RECT 1.410 300.390 3.030 303.870 ;
        RECT 428.830 300.390 430.450 303.870 ;
        RECT 1.410 291.390 3.030 294.870 ;
        RECT 428.830 291.390 430.450 294.870 ;
        RECT 1.410 282.390 3.030 285.870 ;
        RECT 428.830 282.390 430.450 285.870 ;
        RECT 1.410 273.390 3.030 276.870 ;
        RECT 428.830 273.390 430.450 276.870 ;
        RECT 1.410 264.390 3.030 267.870 ;
        RECT 428.830 264.390 430.450 267.870 ;
        RECT 1.410 255.390 3.030 258.870 ;
        RECT 428.830 255.390 430.450 258.870 ;
        RECT 1.410 246.390 3.030 249.870 ;
        RECT 428.830 246.390 430.450 249.870 ;
        RECT 1.410 237.390 3.030 240.870 ;
        RECT 428.830 237.390 430.450 240.870 ;
        RECT 1.410 228.390 3.030 231.870 ;
        RECT 428.830 228.390 430.450 231.870 ;
        RECT 1.410 219.390 3.030 222.870 ;
        RECT 428.830 219.390 430.450 222.870 ;
        RECT 1.410 210.390 3.030 213.870 ;
        RECT 428.830 210.390 430.450 213.870 ;
        RECT 1.410 201.390 3.030 204.870 ;
        RECT 428.830 201.390 430.450 204.870 ;
        RECT 1.410 192.390 3.030 195.870 ;
        RECT 428.830 192.390 430.450 195.870 ;
        RECT 1.410 183.390 3.030 186.870 ;
        RECT 428.830 183.390 430.450 186.870 ;
        RECT 1.410 172.890 3.030 176.370 ;
        RECT 428.830 172.890 430.450 176.370 ;
        RECT 1.410 132.690 3.030 141.750 ;
        RECT 428.830 132.690 430.450 141.750 ;
        RECT 1.410 106.555 3.030 111.275 ;
        RECT 428.830 106.555 430.450 111.275 ;
        RECT 1.410 71.990 3.030 88.490 ;
        RECT 428.830 71.990 430.450 88.490 ;
        RECT 1.410 51.135 3.030 57.095 ;
        RECT 428.830 51.135 430.450 57.095 ;
        RECT 1.410 28.855 3.030 37.915 ;
        RECT 428.830 28.855 430.450 37.915 ;
        RECT 1.410 12.635 3.030 18.595 ;
        RECT 428.830 12.635 430.450 18.595 ;
        RECT 23.210 1.410 28.210 5.000 ;
        RECT 34.635 1.410 35.755 5.000 ;
        RECT 39.730 1.410 40.850 5.000 ;
        RECT 47.210 1.410 52.210 5.000 ;
        RECT 77.210 1.410 82.210 5.000 ;
        RECT 88.635 1.410 89.755 5.000 ;
        RECT 93.730 1.410 94.850 5.000 ;
        RECT 101.210 1.410 106.210 5.000 ;
        RECT 124.280 1.410 125.400 5.000 ;
        RECT 129.365 1.410 130.485 5.000 ;
        RECT 156.620 1.410 161.620 5.000 ;
        RECT 165.110 1.410 170.110 5.000 ;
        RECT 174.155 1.410 179.155 5.000 ;
        RECT 190.140 1.410 195.140 5.000 ;
        RECT 206.165 1.410 211.165 5.000 ;
        RECT 218.165 1.410 223.165 5.000 ;
        RECT 230.165 1.410 235.165 5.000 ;
        RECT 256.165 1.410 261.165 5.000 ;
        RECT 262.390 1.410 267.390 5.000 ;
        RECT 296.565 1.410 297.685 5.000 ;
        RECT 301.650 1.410 302.770 5.000 ;
        RECT 321.090 1.410 326.090 5.000 ;
        RECT 332.515 1.410 333.635 5.000 ;
        RECT 337.610 1.410 338.730 5.000 ;
        RECT 345.090 1.410 350.090 5.000 ;
        RECT 375.090 1.410 380.090 5.000 ;
        RECT 386.515 1.410 387.635 5.000 ;
        RECT 391.610 1.410 392.730 5.000 ;
        RECT 399.090 1.410 404.090 5.000 ;
      LAYER Metal3 ;
        RECT 13.130 481.840 18.130 484.880 ;
        RECT 26.810 481.840 31.810 484.880 ;
        RECT 40.130 481.840 45.130 484.880 ;
        RECT 53.810 481.840 58.810 484.880 ;
        RECT 67.130 481.840 72.130 484.880 ;
        RECT 80.810 481.840 85.810 484.880 ;
        RECT 94.130 481.840 99.130 484.880 ;
        RECT 111.290 481.840 116.290 484.880 ;
        RECT 125.790 481.840 130.790 484.880 ;
        RECT 139.385 481.840 144.385 484.880 ;
        RECT 146.365 481.840 151.365 484.880 ;
        RECT 161.905 481.840 166.905 484.880 ;
        RECT 170.120 481.840 175.120 484.880 ;
        RECT 184.740 481.840 189.740 484.880 ;
        RECT 199.410 481.840 204.410 484.880 ;
        RECT 212.150 481.840 217.150 484.880 ;
        RECT 218.565 481.840 223.565 484.880 ;
        RECT 237.690 481.840 242.690 484.880 ;
        RECT 252.325 481.840 257.325 484.880 ;
        RECT 279.950 481.840 284.950 484.880 ;
        RECT 293.955 481.840 298.955 484.880 ;
        RECT 311.010 481.840 316.010 484.880 ;
        RECT 324.690 481.840 329.690 484.880 ;
        RECT 338.010 481.840 343.010 484.880 ;
        RECT 351.690 481.840 356.690 484.880 ;
        RECT 365.010 481.840 370.010 484.880 ;
        RECT 378.690 481.840 383.690 484.880 ;
        RECT 392.010 481.840 397.010 484.880 ;
        RECT 409.170 481.840 414.170 484.880 ;
        RECT 0.000 471.380 5.000 474.880 ;
        RECT 426.860 471.380 431.860 474.880 ;
        RECT 0.000 462.380 5.000 465.880 ;
        RECT 426.860 462.380 431.860 465.880 ;
        RECT 0.000 453.380 5.000 456.880 ;
        RECT 426.860 453.380 431.860 456.880 ;
        RECT 0.000 444.380 5.000 447.880 ;
        RECT 426.860 444.380 431.860 447.880 ;
        RECT 0.000 435.380 5.000 438.880 ;
        RECT 426.860 435.380 431.860 438.880 ;
        RECT 0.000 426.380 5.000 429.880 ;
        RECT 426.860 426.380 431.860 429.880 ;
        RECT 0.000 417.380 5.000 420.880 ;
        RECT 426.860 417.380 431.860 420.880 ;
        RECT 0.000 408.380 5.000 411.880 ;
        RECT 426.860 408.380 431.860 411.880 ;
        RECT 0.000 399.380 5.000 402.880 ;
        RECT 426.860 399.380 431.860 402.880 ;
        RECT 0.000 390.380 5.000 393.880 ;
        RECT 426.860 390.380 431.860 393.880 ;
        RECT 0.000 381.380 5.000 384.880 ;
        RECT 426.860 381.380 431.860 384.880 ;
        RECT 0.000 372.380 5.000 375.880 ;
        RECT 426.860 372.380 431.860 375.880 ;
        RECT 0.000 363.380 5.000 366.880 ;
        RECT 426.860 363.380 431.860 366.880 ;
        RECT 0.000 354.380 5.000 357.880 ;
        RECT 426.860 354.380 431.860 357.880 ;
        RECT 0.000 345.380 5.000 348.880 ;
        RECT 426.860 345.380 431.860 348.880 ;
        RECT 0.000 336.380 5.000 339.880 ;
        RECT 426.860 336.380 431.860 339.880 ;
        RECT 0.000 327.380 5.000 330.880 ;
        RECT 426.860 327.380 431.860 330.880 ;
        RECT 0.000 318.380 5.000 321.880 ;
        RECT 426.860 318.380 431.860 321.880 ;
        RECT 0.000 309.380 5.000 312.880 ;
        RECT 426.860 309.380 431.860 312.880 ;
        RECT 0.000 300.380 5.000 303.880 ;
        RECT 426.860 300.380 431.860 303.880 ;
        RECT 0.000 291.380 5.000 294.880 ;
        RECT 426.860 291.380 431.860 294.880 ;
        RECT 0.000 282.380 5.000 285.880 ;
        RECT 426.860 282.380 431.860 285.880 ;
        RECT 0.000 273.380 5.000 276.880 ;
        RECT 426.860 273.380 431.860 276.880 ;
        RECT 0.000 264.380 5.000 267.880 ;
        RECT 426.860 264.380 431.860 267.880 ;
        RECT 0.000 255.380 5.000 258.880 ;
        RECT 426.860 255.380 431.860 258.880 ;
        RECT 0.000 246.380 5.000 249.880 ;
        RECT 426.860 246.380 431.860 249.880 ;
        RECT 0.000 237.380 5.000 240.880 ;
        RECT 426.860 237.380 431.860 240.880 ;
        RECT 0.000 228.380 5.000 231.880 ;
        RECT 426.860 228.380 431.860 231.880 ;
        RECT 0.000 219.380 5.000 222.880 ;
        RECT 426.860 219.380 431.860 222.880 ;
        RECT 0.000 210.380 5.000 213.880 ;
        RECT 426.860 210.380 431.860 213.880 ;
        RECT 0.000 201.380 5.000 204.880 ;
        RECT 426.860 201.380 431.860 204.880 ;
        RECT 0.000 192.380 5.000 195.880 ;
        RECT 426.860 192.380 431.860 195.880 ;
        RECT 0.000 183.380 5.000 186.880 ;
        RECT 426.860 183.380 431.860 186.880 ;
        RECT 0.000 172.680 5.000 176.630 ;
        RECT 426.860 172.680 431.860 176.630 ;
        RECT 0.000 132.175 5.000 142.080 ;
        RECT 426.860 132.175 431.860 142.080 ;
        RECT 0.000 106.410 5.000 111.410 ;
        RECT 426.860 106.410 431.860 111.410 ;
        RECT 0.000 71.640 5.000 88.650 ;
        RECT 426.860 71.640 431.860 88.650 ;
        RECT 0.000 50.880 5.000 57.465 ;
        RECT 426.860 50.880 431.860 57.465 ;
        RECT 0.000 28.830 5.000 37.980 ;
        RECT 426.860 28.830 431.860 37.980 ;
        RECT 0.000 12.510 5.000 18.860 ;
        RECT 426.860 12.510 431.860 18.860 ;
        RECT 23.210 0.000 28.210 4.660 ;
        RECT 47.210 0.000 52.210 4.660 ;
        RECT 77.210 0.000 82.210 4.660 ;
        RECT 101.210 0.000 106.210 4.660 ;
        RECT 156.620 0.000 161.620 4.660 ;
        RECT 165.110 0.000 170.110 4.660 ;
        RECT 174.155 0.000 179.155 4.660 ;
        RECT 190.140 0.000 195.140 4.660 ;
        RECT 206.165 0.000 211.165 4.660 ;
        RECT 218.165 0.000 223.165 4.660 ;
        RECT 230.165 0.000 235.165 4.660 ;
        RECT 256.165 0.000 261.165 4.660 ;
        RECT 262.390 0.000 267.390 4.660 ;
        RECT 321.090 0.000 326.090 4.660 ;
        RECT 345.090 0.000 350.090 4.660 ;
        RECT 375.090 0.000 380.090 4.660 ;
        RECT 399.090 0.000 404.090 4.660 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 34.605 132.170 40.815 142.060 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 88.605 132.170 94.815 142.060 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 117.125 132.170 139.140 134.450 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.245 50.870 121.250 57.455 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126.880 472.305 129.740 473.925 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.010 472.630 273.110 473.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.275 472.305 297.135 473.925 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 463.630 273.110 464.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 454.630 273.110 455.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 445.630 273.110 446.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 436.630 273.110 437.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 427.630 273.110 428.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 418.630 273.110 419.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 409.630 273.110 410.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 400.630 273.110 401.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 391.630 273.110 392.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 382.630 273.110 383.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 373.630 273.110 374.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 364.630 273.110 365.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 355.630 273.110 356.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 346.630 273.110 347.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 337.630 273.110 338.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 328.630 273.110 329.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 319.630 273.110 320.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 310.630 273.110 311.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 301.630 273.110 302.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 292.630 273.110 293.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 283.630 273.110 284.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 274.630 273.110 275.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 265.630 273.110 266.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 256.630 273.110 257.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 247.630 273.110 248.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 238.630 273.110 239.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 229.630 273.110 230.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 220.630 273.110 221.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 211.630 273.110 212.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 202.630 273.110 203.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 193.630 273.110 194.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 152.015 184.630 273.110 185.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 332.485 132.170 338.695 142.060 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 386.485 132.170 392.695 142.060 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.180 109.130 139.130 111.410 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 280.390 109.130 288.405 115.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 120.555 71.645 139.140 82.990 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.390 66.215 229.885 75.075 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.475 71.635 418.815 83.920 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 50.865 422.410 57.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 11.245 34.900 121.250 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.435 30.885 206.985 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.565 39.500 206.985 42.910 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 174.300 32.960 277.410 36.960 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 209.285 45.825 257.150 52.100 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.610 28.830 312.145 30.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 309.125 34.900 423.935 37.975 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 137.190 17.620 138.890 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 143.820 17.620 144.470 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 208.870 17.620 209.520 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 211.495 17.620 212.145 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 234.365 17.620 235.015 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 236.605 17.620 237.255 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 238.845 17.620 239.495 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 241.085 17.620 241.735 19.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.725 17.620 306.075 19.380 ;
    END
  END VSS
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 413.475 0.000 414.595 5.000 ;
    END
  END WEN[7]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 363.150 0.000 364.270 5.000 ;
    END
  END WEN[6]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 360.900 0.000 362.020 5.000 ;
    END
  END WEN[5]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 310.575 0.000 311.695 5.000 ;
    END
  END WEN[4]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.020 0.000 118.140 5.000 ;
    END
  END WEN[3]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.270 0.000 66.390 5.000 ;
    END
  END WEN[2]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.020 0.000 64.140 5.000 ;
    END
  END WEN[1]
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.938000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.695 0.000 13.815 5.000 ;
    END
  END WEN[0]
  OBS
      LAYER Metal1 ;
        RECT 5.000 5.000 426.860 479.880 ;
      LAYER Metal2 ;
        RECT 5.000 5.000 426.860 479.880 ;
      LAYER Metal3 ;
        RECT 5.000 5.000 426.860 479.880 ;
  END
END gf180mcu_fd_ip_sram__sram512x8m8wm1
END LIBRARY

