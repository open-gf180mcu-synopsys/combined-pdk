magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1900 1270
<< nmos >>
rect 200 210 260 380
rect 400 210 460 380
rect 540 210 600 380
rect 710 210 770 380
rect 950 210 1010 380
rect 1150 210 1210 380
rect 1470 210 1530 380
rect 1640 210 1700 380
<< pmos >>
rect 200 720 260 1060
rect 370 720 430 1060
rect 540 720 600 1060
rect 710 720 770 1060
rect 980 720 1040 1060
rect 1150 720 1210 1060
rect 1470 720 1530 1060
rect 1640 720 1700 1060
<< ndiff >>
rect 100 318 200 380
rect 100 272 122 318
rect 168 272 200 318
rect 100 210 200 272
rect 260 288 400 380
rect 260 242 307 288
rect 353 242 400 288
rect 260 210 400 242
rect 460 210 540 380
rect 600 293 710 380
rect 600 247 632 293
rect 678 247 710 293
rect 600 210 710 247
rect 770 210 950 380
rect 1010 283 1150 380
rect 1010 237 1057 283
rect 1103 237 1150 283
rect 1010 210 1150 237
rect 1210 318 1310 380
rect 1210 272 1242 318
rect 1288 272 1310 318
rect 1210 210 1310 272
rect 1370 318 1470 380
rect 1370 272 1392 318
rect 1438 272 1470 318
rect 1370 210 1470 272
rect 1530 283 1640 380
rect 1530 237 1562 283
rect 1608 237 1640 283
rect 1530 210 1640 237
rect 1700 318 1800 380
rect 1700 272 1732 318
rect 1778 272 1800 318
rect 1700 210 1800 272
<< pdiff >>
rect 100 1007 200 1060
rect 100 773 122 1007
rect 168 773 200 1007
rect 100 720 200 773
rect 260 1040 370 1060
rect 260 900 292 1040
rect 338 900 370 1040
rect 260 720 370 900
rect 430 720 540 1060
rect 600 1037 710 1060
rect 600 803 632 1037
rect 678 803 710 1037
rect 600 720 710 803
rect 770 720 980 1060
rect 1040 1032 1150 1060
rect 1040 798 1072 1032
rect 1118 798 1150 1032
rect 1040 720 1150 798
rect 1210 1037 1310 1060
rect 1210 803 1242 1037
rect 1288 803 1310 1037
rect 1210 720 1310 803
rect 1370 1012 1470 1060
rect 1370 778 1392 1012
rect 1438 778 1470 1012
rect 1370 720 1470 778
rect 1530 1030 1640 1060
rect 1530 890 1562 1030
rect 1608 890 1640 1030
rect 1530 720 1640 890
rect 1700 1007 1800 1060
rect 1700 773 1732 1007
rect 1778 773 1800 1007
rect 1700 720 1800 773
<< ndiffc >>
rect 122 272 168 318
rect 307 242 353 288
rect 632 247 678 293
rect 1057 237 1103 283
rect 1242 272 1288 318
rect 1392 272 1438 318
rect 1562 237 1608 283
rect 1732 272 1778 318
<< pdiffc >>
rect 122 773 168 1007
rect 292 900 338 1040
rect 632 803 678 1037
rect 1072 798 1118 1032
rect 1242 803 1288 1037
rect 1392 778 1438 1012
rect 1562 890 1608 1030
rect 1732 773 1778 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 310 118 460 140
rect 310 72 362 118
rect 408 72 460 118
rect 310 50 460 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1030 118 1180 140
rect 1030 72 1082 118
rect 1128 72 1180 118
rect 1030 50 1180 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 310 1198 460 1220
rect 310 1152 362 1198
rect 408 1152 460 1198
rect 310 1130 460 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1030 1198 1180 1220
rect 1030 1152 1082 1198
rect 1128 1152 1180 1198
rect 1030 1130 1180 1152
rect 1270 1198 1420 1220
rect 1270 1152 1322 1198
rect 1368 1152 1420 1198
rect 1270 1130 1420 1152
rect 1510 1198 1660 1220
rect 1510 1152 1562 1198
rect 1608 1152 1660 1198
rect 1510 1130 1660 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 362 72 408 118
rect 592 72 638 118
rect 832 72 878 118
rect 1082 72 1128 118
rect 1312 72 1358 118
rect 1552 72 1598 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 362 1152 408 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1082 1152 1128 1198
rect 1322 1152 1368 1198
rect 1562 1152 1608 1198
<< polysilicon >>
rect 200 1060 260 1110
rect 370 1060 430 1110
rect 540 1060 600 1110
rect 710 1060 770 1110
rect 980 1060 1040 1110
rect 1150 1060 1210 1110
rect 1470 1060 1530 1110
rect 1640 1060 1700 1110
rect 200 700 260 720
rect 200 673 320 700
rect 200 627 237 673
rect 283 627 320 673
rect 200 600 320 627
rect 370 670 430 720
rect 540 700 600 720
rect 710 700 770 720
rect 520 673 620 700
rect 370 643 470 670
rect 200 380 260 600
rect 370 597 397 643
rect 443 597 470 643
rect 520 627 547 673
rect 593 627 620 673
rect 520 600 620 627
rect 680 673 780 700
rect 680 627 707 673
rect 753 627 780 673
rect 680 600 780 627
rect 370 570 470 597
rect 370 440 430 570
rect 710 550 770 600
rect 540 510 770 550
rect 830 563 930 590
rect 830 517 857 563
rect 903 517 930 563
rect 370 400 460 440
rect 400 380 460 400
rect 540 380 600 510
rect 830 490 930 517
rect 980 570 1040 720
rect 1150 700 1210 720
rect 1140 673 1240 700
rect 1140 627 1167 673
rect 1213 627 1240 673
rect 1140 600 1240 627
rect 980 543 1100 570
rect 980 497 1027 543
rect 1073 497 1100 543
rect 830 460 900 490
rect 710 420 900 460
rect 980 470 1100 497
rect 980 440 1040 470
rect 710 380 770 420
rect 950 400 1040 440
rect 950 380 1010 400
rect 1150 380 1210 600
rect 1470 570 1530 720
rect 1640 570 1700 720
rect 1440 548 1530 570
rect 1440 502 1462 548
rect 1508 502 1530 548
rect 1440 480 1530 502
rect 1470 380 1530 480
rect 1580 543 1700 570
rect 1580 497 1607 543
rect 1653 497 1700 543
rect 1580 470 1700 497
rect 1640 380 1700 470
rect 200 160 260 210
rect 400 160 460 210
rect 540 160 600 210
rect 710 160 770 210
rect 950 160 1010 210
rect 1150 160 1210 210
rect 1470 160 1530 210
rect 1640 160 1700 210
<< polycontact >>
rect 237 627 283 673
rect 397 597 443 643
rect 547 627 593 673
rect 707 627 753 673
rect 857 517 903 563
rect 1167 627 1213 673
rect 1027 497 1073 543
rect 1462 502 1508 548
rect 1607 497 1653 543
<< metal1 >>
rect 0 1198 1900 1270
rect 0 1152 112 1198
rect 158 1152 362 1198
rect 408 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1082 1198
rect 1128 1152 1322 1198
rect 1368 1152 1562 1198
rect 1608 1152 1900 1198
rect 0 1130 1900 1152
rect 120 1007 170 1060
rect 120 773 122 1007
rect 168 773 170 1007
rect 290 1040 340 1130
rect 290 900 292 1040
rect 338 900 340 1040
rect 290 880 340 900
rect 630 1037 680 1060
rect 630 830 632 1037
rect 120 530 170 773
rect 230 803 632 830
rect 678 803 680 1037
rect 230 780 680 803
rect 1070 1032 1120 1130
rect 1070 798 1072 1032
rect 1118 798 1120 1032
rect 230 680 280 780
rect 1070 770 1120 798
rect 1240 1037 1290 1060
rect 1240 803 1242 1037
rect 1288 803 1290 1037
rect 1240 800 1290 803
rect 1390 1012 1440 1060
rect 1240 750 1340 800
rect 220 673 310 680
rect 220 627 237 673
rect 283 627 310 673
rect 520 673 620 680
rect 220 620 310 627
rect 370 646 470 650
rect 100 520 170 530
rect 70 516 170 520
rect 70 464 94 516
rect 146 464 170 516
rect 70 460 170 464
rect 90 450 170 460
rect 120 318 170 450
rect 230 450 280 620
rect 370 594 394 646
rect 446 594 470 646
rect 520 627 547 673
rect 593 627 620 673
rect 520 620 620 627
rect 680 673 780 680
rect 680 646 707 673
rect 753 646 780 673
rect 370 590 470 594
rect 540 540 600 620
rect 680 594 704 646
rect 756 594 780 646
rect 1140 676 1240 680
rect 1140 624 1164 676
rect 1216 624 1240 676
rect 1140 620 1240 624
rect 680 590 780 594
rect 830 563 930 570
rect 830 540 857 563
rect 540 517 857 540
rect 903 517 930 563
rect 540 510 930 517
rect 1000 546 1100 550
rect 540 490 910 510
rect 1000 494 1024 546
rect 1076 494 1100 546
rect 1000 490 1100 494
rect 540 480 900 490
rect 230 400 480 450
rect 120 272 122 318
rect 168 272 170 318
rect 120 210 170 272
rect 290 288 370 320
rect 290 242 307 288
rect 353 242 370 288
rect 430 310 480 400
rect 840 410 900 480
rect 1290 470 1340 750
rect 1390 778 1392 1012
rect 1438 778 1440 1012
rect 1560 1030 1610 1130
rect 1560 890 1562 1030
rect 1608 890 1610 1030
rect 1560 860 1610 890
rect 1730 1007 1780 1060
rect 1390 740 1440 778
rect 1730 773 1732 1007
rect 1778 773 1780 1007
rect 1390 690 1660 740
rect 1440 548 1540 550
rect 1440 502 1462 548
rect 1508 546 1540 548
rect 1440 494 1464 502
rect 1516 494 1540 546
rect 1440 490 1540 494
rect 1600 543 1660 690
rect 1600 497 1607 543
rect 1653 497 1660 543
rect 1240 420 1340 470
rect 1600 440 1660 497
rect 1240 410 1290 420
rect 840 360 1290 410
rect 630 310 680 330
rect 1240 318 1290 360
rect 430 293 680 310
rect 430 260 632 293
rect 290 140 370 242
rect 630 247 632 260
rect 678 247 680 293
rect 630 210 680 247
rect 1040 283 1120 310
rect 1040 237 1057 283
rect 1103 237 1120 283
rect 1040 140 1120 237
rect 1240 272 1242 318
rect 1288 272 1290 318
rect 1240 210 1290 272
rect 1390 390 1660 440
rect 1730 660 1780 773
rect 1730 650 1810 660
rect 1730 646 1830 650
rect 1730 594 1754 646
rect 1806 594 1830 646
rect 1730 590 1830 594
rect 1730 580 1810 590
rect 1390 318 1440 390
rect 1390 272 1392 318
rect 1438 272 1440 318
rect 1730 318 1780 580
rect 1390 210 1440 272
rect 1560 283 1610 310
rect 1560 237 1562 283
rect 1608 237 1610 283
rect 1560 140 1610 237
rect 1730 272 1732 318
rect 1778 272 1780 318
rect 1730 210 1780 272
rect 0 118 1900 140
rect 0 72 112 118
rect 158 72 362 118
rect 408 72 592 118
rect 638 72 832 118
rect 878 72 1082 118
rect 1128 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1900 118
rect 0 0 1900 72
<< via1 >>
rect 94 464 146 516
rect 394 643 446 646
rect 394 597 397 643
rect 397 597 443 643
rect 443 597 446 643
rect 394 594 446 597
rect 704 627 707 646
rect 707 627 753 646
rect 753 627 756 646
rect 704 594 756 627
rect 1164 673 1216 676
rect 1164 627 1167 673
rect 1167 627 1213 673
rect 1213 627 1216 673
rect 1164 624 1216 627
rect 1024 543 1076 546
rect 1024 497 1027 543
rect 1027 497 1073 543
rect 1073 497 1076 543
rect 1024 494 1076 497
rect 1464 502 1508 546
rect 1508 502 1516 546
rect 1464 494 1516 502
rect 1754 594 1806 646
<< metal2 >>
rect 1140 680 1240 690
rect 700 676 1240 680
rect 700 660 1164 676
rect 370 646 470 660
rect 690 650 1164 660
rect 370 594 394 646
rect 446 594 470 646
rect 370 580 470 594
rect 680 646 1164 650
rect 680 594 704 646
rect 756 624 1164 646
rect 1216 624 1240 676
rect 1740 650 1820 660
rect 756 620 1240 624
rect 756 594 780 620
rect 1140 610 1240 620
rect 1730 646 1830 650
rect 680 590 780 594
rect 1730 594 1754 646
rect 1806 594 1830 646
rect 1730 590 1830 594
rect 690 580 770 590
rect 1740 580 1820 590
rect 1010 550 1090 560
rect 1440 550 1540 560
rect 920 546 1540 550
rect 70 520 170 530
rect 920 520 1024 546
rect 70 516 1024 520
rect 70 464 94 516
rect 146 494 1024 516
rect 1076 494 1464 546
rect 1516 494 1540 546
rect 146 490 1540 494
rect 146 480 1090 490
rect 1440 480 1540 490
rect 146 464 980 480
rect 70 460 980 464
rect 70 450 170 460
<< labels >>
rlabel via1 s 394 594 446 646 4 D
port 1 nsew signal input
rlabel via1 s 1754 594 1806 646 4 Q
port 2 nsew signal output
rlabel via1 s 1164 624 1216 676 4 CLK
port 3 nsew clock input
rlabel metal1 s 290 880 340 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 0 370 320 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1070 770 1120 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1560 860 1610 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1900 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1040 0 1120 310 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1560 0 1610 310 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1900 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 704 594 756 646 1 CLK
port 3 nsew clock input
rlabel metal2 s 690 580 770 660 1 CLK
port 3 nsew clock input
rlabel metal2 s 680 590 780 650 1 CLK
port 3 nsew clock input
rlabel metal2 s 700 620 1240 680 1 CLK
port 3 nsew clock input
rlabel metal2 s 1140 610 1240 690 1 CLK
port 3 nsew clock input
rlabel metal1 s 680 590 780 680 1 CLK
port 3 nsew clock input
rlabel metal1 s 1140 620 1240 680 1 CLK
port 3 nsew clock input
rlabel metal2 s 370 580 470 660 1 D
port 1 nsew signal input
rlabel metal1 s 370 590 470 650 1 D
port 1 nsew signal input
rlabel metal2 s 1740 580 1820 660 1 Q
port 2 nsew signal output
rlabel metal2 s 1730 590 1830 650 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 210 1780 1060 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 580 1810 660 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 590 1830 650 1 Q
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1900 1270
string GDS_END 266016
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 252440
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
