magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 780 1270
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
rect 500 210 560 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
<< ndiff >>
rect 120 318 220 380
rect 120 272 142 318
rect 188 272 220 318
rect 120 210 220 272
rect 280 210 330 380
rect 390 303 500 380
rect 390 257 422 303
rect 468 257 500 303
rect 390 210 500 257
rect 560 278 660 380
rect 560 232 592 278
rect 638 232 660 278
rect 560 210 660 232
<< pdiff >>
rect 90 1035 190 1060
rect 90 895 112 1035
rect 158 895 190 1035
rect 90 720 190 895
rect 250 1035 360 1060
rect 250 895 282 1035
rect 328 895 360 1035
rect 250 720 360 895
rect 420 1035 530 1060
rect 420 895 452 1035
rect 498 895 530 1035
rect 420 720 530 895
rect 590 1040 690 1060
rect 590 900 622 1040
rect 668 900 690 1040
rect 590 720 690 900
<< ndiffc >>
rect 142 272 188 318
rect 422 257 468 303
rect 592 232 638 278
<< pdiffc >>
rect 112 895 158 1035
rect 282 895 328 1035
rect 452 895 498 1035
rect 622 900 668 1040
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 190 540 250 720
rect 360 670 420 720
rect 300 643 420 670
rect 300 597 347 643
rect 393 597 420 643
rect 300 570 420 597
rect 110 513 250 540
rect 110 467 147 513
rect 193 467 250 513
rect 110 450 250 467
rect 360 450 420 570
rect 530 540 590 720
rect 110 440 280 450
rect 190 410 280 440
rect 220 380 280 410
rect 330 400 420 450
rect 470 513 590 540
rect 470 467 497 513
rect 543 467 590 513
rect 470 440 590 467
rect 330 380 390 400
rect 500 380 560 440
rect 220 160 280 210
rect 330 160 390 210
rect 500 160 560 210
<< polycontact >>
rect 347 597 393 643
rect 147 467 193 513
rect 497 467 543 513
<< metal1 >>
rect 0 1198 780 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 780 1198
rect 0 1130 780 1152
rect 110 1035 160 1060
rect 110 895 112 1035
rect 158 895 160 1035
rect 110 820 160 895
rect 280 1035 330 1130
rect 280 895 282 1035
rect 328 895 330 1035
rect 280 870 330 895
rect 450 1035 500 1060
rect 450 895 452 1035
rect 498 895 500 1035
rect 450 820 500 895
rect 110 770 500 820
rect 620 1040 670 1060
rect 620 900 622 1040
rect 668 900 670 1040
rect 620 780 670 900
rect 600 776 700 780
rect 600 724 624 776
rect 676 724 700 776
rect 600 720 700 724
rect 320 646 420 650
rect 320 594 344 646
rect 396 594 420 646
rect 320 590 420 594
rect 120 516 220 520
rect 120 464 144 516
rect 196 464 220 516
rect 120 460 220 464
rect 470 516 570 520
rect 470 464 494 516
rect 546 464 570 516
rect 470 460 570 464
rect 620 400 670 720
rect 140 318 190 380
rect 140 272 142 318
rect 188 272 190 318
rect 140 140 190 272
rect 420 350 670 400
rect 420 303 470 350
rect 420 257 422 303
rect 468 257 470 303
rect 420 210 470 257
rect 590 278 640 300
rect 590 232 592 278
rect 638 232 640 278
rect 590 140 640 232
rect 0 118 780 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 780 118
rect 0 0 780 72
<< via1 >>
rect 624 724 676 776
rect 344 643 396 646
rect 344 597 347 643
rect 347 597 393 643
rect 393 597 396 643
rect 344 594 396 597
rect 144 513 196 516
rect 144 467 147 513
rect 147 467 193 513
rect 193 467 196 513
rect 144 464 196 467
rect 494 513 546 516
rect 494 467 497 513
rect 497 467 543 513
rect 543 467 546 513
rect 494 464 546 467
<< metal2 >>
rect 600 776 700 790
rect 600 724 624 776
rect 676 724 700 776
rect 600 710 700 724
rect 320 646 420 660
rect 320 594 344 646
rect 396 594 420 646
rect 320 580 420 594
rect 120 516 220 530
rect 120 464 144 516
rect 196 464 220 516
rect 120 450 220 464
rect 470 516 570 530
rect 470 464 494 516
rect 546 464 570 516
rect 470 450 570 464
<< labels >>
rlabel via1 s 624 724 676 776 4 Y
port 1 nsew signal output
rlabel via1 s 144 464 196 516 4 A0
port 2 nsew signal input
rlabel via1 s 344 594 396 646 4 A1
port 3 nsew signal input
rlabel via1 s 494 464 546 516 4 B
port 4 nsew signal input
rlabel metal1 s 280 870 330 1270 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 140 0 190 380 4 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 1130 780 1270 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 590 0 640 300 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 0 780 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal2 s 120 450 220 530 1 A0
port 2 nsew signal input
rlabel metal1 s 120 460 220 520 1 A0
port 2 nsew signal input
rlabel metal2 s 320 580 420 660 1 A1
port 3 nsew signal input
rlabel metal1 s 320 590 420 650 1 A1
port 3 nsew signal input
rlabel metal2 s 470 450 570 530 1 B
port 4 nsew signal input
rlabel metal1 s 470 460 570 520 1 B
port 4 nsew signal input
rlabel metal2 s 600 710 700 790 1 Y
port 1 nsew signal output
rlabel metal1 s 420 210 470 400 1 Y
port 1 nsew signal output
rlabel metal1 s 420 350 670 400 1 Y
port 1 nsew signal output
rlabel metal1 s 620 350 670 1060 1 Y
port 1 nsew signal output
rlabel metal1 s 600 720 700 780 1 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 780 1270
string GDS_END 46002
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 40774
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
