magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 760 220 830
rect 55 555 80 760
rect 140 520 165 725
rect 130 518 180 520
rect 130 492 142 518
rect 168 492 180 518
rect 130 490 180 492
rect 140 485 165 490
rect 55 70 80 190
rect 0 0 220 70
<< via1 >>
rect 142 492 168 518
<< obsm1 >>
rect 115 230 165 255
rect 140 105 165 230
<< metal2 >>
rect 130 518 180 525
rect 130 492 142 518
rect 168 492 180 518
rect 130 485 180 492
<< labels >>
rlabel metal1 s 55 555 80 830 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 760 220 830 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 55 0 80 190 6 VSS
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 0 220 70 6 VSS
port 3 nsew ground bidirectional abutment
rlabel via1 s 142 492 168 518 6 Y
port 1 nsew signal output
rlabel metal2 s 130 485 180 525 6 Y
port 1 nsew signal output
rlabel metal1 s 140 485 165 725 6 Y
port 1 nsew signal output
rlabel metal1 s 130 490 180 520 6 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 220 830
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 507132
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 504578
<< end >>
