magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 3160 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 530 210 590 380
rect 700 210 760 380
rect 870 210 930 380
rect 1040 210 1100 380
rect 1210 210 1270 380
rect 1380 210 1440 380
rect 1550 210 1610 380
rect 1720 210 1780 380
rect 1890 210 1950 380
rect 2060 210 2120 380
rect 2230 210 2290 380
rect 2400 210 2460 380
rect 2570 210 2630 380
rect 2740 210 2800 380
rect 2910 210 2970 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
rect 700 720 760 1060
rect 870 720 930 1060
rect 1040 720 1100 1060
rect 1210 720 1270 1060
rect 1380 720 1440 1060
rect 1550 720 1610 1060
rect 1720 720 1780 1060
rect 1890 720 1950 1060
rect 2060 720 2120 1060
rect 2230 720 2290 1060
rect 2400 720 2460 1060
rect 2570 720 2630 1060
rect 2740 720 2800 1060
rect 2910 720 2970 1060
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 318 530 380
rect 420 272 452 318
rect 498 272 530 318
rect 420 210 530 272
rect 590 318 700 380
rect 590 272 622 318
rect 668 272 700 318
rect 590 210 700 272
rect 760 318 870 380
rect 760 272 792 318
rect 838 272 870 318
rect 760 210 870 272
rect 930 318 1040 380
rect 930 272 962 318
rect 1008 272 1040 318
rect 930 210 1040 272
rect 1100 318 1210 380
rect 1100 272 1132 318
rect 1178 272 1210 318
rect 1100 210 1210 272
rect 1270 318 1380 380
rect 1270 272 1302 318
rect 1348 272 1380 318
rect 1270 210 1380 272
rect 1440 318 1550 380
rect 1440 272 1472 318
rect 1518 272 1550 318
rect 1440 210 1550 272
rect 1610 318 1720 380
rect 1610 272 1642 318
rect 1688 272 1720 318
rect 1610 210 1720 272
rect 1780 318 1890 380
rect 1780 272 1812 318
rect 1858 272 1890 318
rect 1780 210 1890 272
rect 1950 318 2060 380
rect 1950 272 1982 318
rect 2028 272 2060 318
rect 1950 210 2060 272
rect 2120 318 2230 380
rect 2120 272 2152 318
rect 2198 272 2230 318
rect 2120 210 2230 272
rect 2290 318 2400 380
rect 2290 272 2322 318
rect 2368 272 2400 318
rect 2290 210 2400 272
rect 2460 318 2570 380
rect 2460 272 2492 318
rect 2538 272 2570 318
rect 2460 210 2570 272
rect 2630 318 2740 380
rect 2630 272 2662 318
rect 2708 272 2740 318
rect 2630 210 2740 272
rect 2800 318 2910 380
rect 2800 272 2832 318
rect 2878 272 2910 318
rect 2800 210 2910 272
rect 2970 318 3070 380
rect 2970 272 3002 318
rect 3048 272 3070 318
rect 2970 210 3070 272
<< pdiff >>
rect 90 1007 190 1060
rect 90 773 112 1007
rect 158 773 190 1007
rect 90 720 190 773
rect 250 1007 360 1060
rect 250 773 282 1007
rect 328 773 360 1007
rect 250 720 360 773
rect 420 1032 530 1060
rect 420 798 452 1032
rect 498 798 530 1032
rect 420 720 530 798
rect 590 1007 700 1060
rect 590 773 622 1007
rect 668 773 700 1007
rect 590 720 700 773
rect 760 1032 870 1060
rect 760 798 792 1032
rect 838 798 870 1032
rect 760 720 870 798
rect 930 1007 1040 1060
rect 930 773 962 1007
rect 1008 773 1040 1007
rect 930 720 1040 773
rect 1100 1032 1210 1060
rect 1100 798 1132 1032
rect 1178 798 1210 1032
rect 1100 720 1210 798
rect 1270 1007 1380 1060
rect 1270 773 1302 1007
rect 1348 773 1380 1007
rect 1270 720 1380 773
rect 1440 1032 1550 1060
rect 1440 798 1472 1032
rect 1518 798 1550 1032
rect 1440 720 1550 798
rect 1610 1007 1720 1060
rect 1610 773 1642 1007
rect 1688 773 1720 1007
rect 1610 720 1720 773
rect 1780 1032 1890 1060
rect 1780 798 1812 1032
rect 1858 798 1890 1032
rect 1780 720 1890 798
rect 1950 1007 2060 1060
rect 1950 773 1982 1007
rect 2028 773 2060 1007
rect 1950 720 2060 773
rect 2120 1032 2230 1060
rect 2120 798 2152 1032
rect 2198 798 2230 1032
rect 2120 720 2230 798
rect 2290 1007 2400 1060
rect 2290 773 2322 1007
rect 2368 773 2400 1007
rect 2290 720 2400 773
rect 2460 1032 2570 1060
rect 2460 798 2492 1032
rect 2538 798 2570 1032
rect 2460 720 2570 798
rect 2630 1007 2740 1060
rect 2630 773 2662 1007
rect 2708 773 2740 1007
rect 2630 720 2740 773
rect 2800 1032 2910 1060
rect 2800 798 2832 1032
rect 2878 798 2910 1032
rect 2800 720 2910 798
rect 2970 1007 3070 1060
rect 2970 773 3002 1007
rect 3048 773 3070 1007
rect 2970 720 3070 773
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 792 272 838 318
rect 962 272 1008 318
rect 1132 272 1178 318
rect 1302 272 1348 318
rect 1472 272 1518 318
rect 1642 272 1688 318
rect 1812 272 1858 318
rect 1982 272 2028 318
rect 2152 272 2198 318
rect 2322 272 2368 318
rect 2492 272 2538 318
rect 2662 272 2708 318
rect 2832 272 2878 318
rect 3002 272 3048 318
<< pdiffc >>
rect 112 773 158 1007
rect 282 773 328 1007
rect 452 798 498 1032
rect 622 773 668 1007
rect 792 798 838 1032
rect 962 773 1008 1007
rect 1132 798 1178 1032
rect 1302 773 1348 1007
rect 1472 798 1518 1032
rect 1642 773 1688 1007
rect 1812 798 1858 1032
rect 1982 773 2028 1007
rect 2152 798 2198 1032
rect 2322 773 2368 1007
rect 2492 798 2538 1032
rect 2662 773 2708 1007
rect 2832 798 2878 1032
rect 3002 773 3048 1007
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
rect 1260 118 1410 140
rect 1260 72 1312 118
rect 1358 72 1410 118
rect 1260 50 1410 72
rect 1500 118 1650 140
rect 1500 72 1552 118
rect 1598 72 1650 118
rect 1500 50 1650 72
rect 1740 118 1890 140
rect 1740 72 1792 118
rect 1838 72 1890 118
rect 1740 50 1890 72
rect 1980 118 2130 140
rect 1980 72 2032 118
rect 2078 72 2130 118
rect 1980 50 2130 72
rect 2220 118 2370 140
rect 2220 72 2272 118
rect 2318 72 2370 118
rect 2220 50 2370 72
rect 2460 118 2610 140
rect 2460 72 2512 118
rect 2558 72 2610 118
rect 2460 50 2610 72
rect 2700 118 2850 140
rect 2700 72 2752 118
rect 2798 72 2850 118
rect 2700 50 2850 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
rect 1260 1198 1410 1220
rect 1260 1152 1312 1198
rect 1358 1152 1410 1198
rect 1260 1130 1410 1152
rect 1500 1198 1650 1220
rect 1500 1152 1552 1198
rect 1598 1152 1650 1198
rect 1500 1130 1650 1152
rect 1740 1198 1890 1220
rect 1740 1152 1792 1198
rect 1838 1152 1890 1198
rect 1740 1130 1890 1152
rect 1980 1198 2130 1220
rect 1980 1152 2032 1198
rect 2078 1152 2130 1198
rect 1980 1130 2130 1152
rect 2220 1198 2370 1220
rect 2220 1152 2272 1198
rect 2318 1152 2370 1198
rect 2220 1130 2370 1152
rect 2460 1198 2610 1220
rect 2460 1152 2512 1198
rect 2558 1152 2610 1198
rect 2460 1130 2610 1152
rect 2700 1198 2850 1220
rect 2700 1152 2752 1198
rect 2798 1152 2850 1198
rect 2700 1130 2850 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
rect 1312 72 1358 118
rect 1552 72 1598 118
rect 1792 72 1838 118
rect 2032 72 2078 118
rect 2272 72 2318 118
rect 2512 72 2558 118
rect 2752 72 2798 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
rect 1312 1152 1358 1198
rect 1552 1152 1598 1198
rect 1792 1152 1838 1198
rect 2032 1152 2078 1198
rect 2272 1152 2318 1198
rect 2512 1152 2558 1198
rect 2752 1152 2798 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 700 1060 760 1110
rect 870 1060 930 1110
rect 1040 1060 1100 1110
rect 1210 1060 1270 1110
rect 1380 1060 1440 1110
rect 1550 1060 1610 1110
rect 1720 1060 1780 1110
rect 1890 1060 1950 1110
rect 2060 1060 2120 1110
rect 2230 1060 2290 1110
rect 2400 1060 2460 1110
rect 2570 1060 2630 1110
rect 2740 1060 2800 1110
rect 2910 1060 2970 1110
rect 190 540 250 720
rect 360 700 420 720
rect 530 700 590 720
rect 700 700 760 720
rect 870 700 930 720
rect 1040 700 1100 720
rect 1210 700 1270 720
rect 1380 700 1440 720
rect 1550 700 1610 720
rect 1720 700 1780 720
rect 1890 700 1950 720
rect 2060 700 2120 720
rect 2230 700 2290 720
rect 2400 700 2460 720
rect 2570 700 2630 720
rect 2740 700 2800 720
rect 2910 700 2970 720
rect 360 690 2970 700
rect 300 663 2970 690
rect 300 617 327 663
rect 373 640 2970 663
rect 373 617 420 640
rect 300 590 420 617
rect 190 513 310 540
rect 190 467 237 513
rect 283 467 310 513
rect 190 440 310 467
rect 360 460 420 590
rect 700 460 760 640
rect 1040 460 1100 640
rect 1380 460 1440 640
rect 1720 460 1780 640
rect 2060 460 2120 640
rect 2400 460 2460 640
rect 2740 460 2800 640
rect 190 380 250 440
rect 360 400 2970 460
rect 360 380 420 400
rect 530 380 590 400
rect 700 380 760 400
rect 870 380 930 400
rect 1040 380 1100 400
rect 1210 380 1270 400
rect 1380 380 1440 400
rect 1550 380 1610 400
rect 1720 380 1780 400
rect 1890 380 1950 400
rect 2060 380 2120 400
rect 2230 380 2290 400
rect 2400 380 2460 400
rect 2570 380 2630 400
rect 2740 380 2800 400
rect 2910 380 2970 400
rect 190 160 250 210
rect 360 160 420 210
rect 530 160 590 210
rect 700 160 760 210
rect 870 160 930 210
rect 1040 160 1100 210
rect 1210 160 1270 210
rect 1380 160 1440 210
rect 1550 160 1610 210
rect 1720 160 1780 210
rect 1890 160 1950 210
rect 2060 160 2120 210
rect 2230 160 2290 210
rect 2400 160 2460 210
rect 2570 160 2630 210
rect 2740 160 2800 210
rect 2910 160 2970 210
<< polycontact >>
rect 327 617 373 663
rect 237 467 283 513
<< metal1 >>
rect 0 1198 3160 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1312 1198
rect 1358 1152 1552 1198
rect 1598 1152 1792 1198
rect 1838 1152 2032 1198
rect 2078 1152 2272 1198
rect 2318 1152 2512 1198
rect 2558 1152 2752 1198
rect 2798 1152 3160 1198
rect 0 1130 3160 1152
rect 110 1007 160 1060
rect 110 773 112 1007
rect 158 773 160 1007
rect 110 670 160 773
rect 280 1007 330 1130
rect 280 773 282 1007
rect 328 773 330 1007
rect 280 720 330 773
rect 450 1032 500 1060
rect 450 798 452 1032
rect 498 798 500 1032
rect 450 670 500 798
rect 620 1007 670 1130
rect 620 773 622 1007
rect 668 773 670 1007
rect 620 720 670 773
rect 790 1032 840 1060
rect 790 798 792 1032
rect 838 798 840 1032
rect 790 670 840 798
rect 960 1007 1010 1130
rect 960 773 962 1007
rect 1008 773 1010 1007
rect 960 720 1010 773
rect 1130 1032 1180 1060
rect 1130 798 1132 1032
rect 1178 798 1180 1032
rect 1130 670 1180 798
rect 1300 1007 1350 1130
rect 1300 773 1302 1007
rect 1348 773 1350 1007
rect 1300 720 1350 773
rect 1470 1032 1520 1060
rect 1470 798 1472 1032
rect 1518 798 1520 1032
rect 1470 670 1520 798
rect 1640 1007 1690 1130
rect 1640 773 1642 1007
rect 1688 773 1690 1007
rect 1640 720 1690 773
rect 1810 1032 1860 1060
rect 1810 798 1812 1032
rect 1858 798 1860 1032
rect 1810 670 1860 798
rect 1980 1007 2030 1130
rect 1980 773 1982 1007
rect 2028 773 2030 1007
rect 1980 720 2030 773
rect 2150 1032 2200 1060
rect 2150 798 2152 1032
rect 2198 798 2200 1032
rect 2150 670 2200 798
rect 2320 1007 2370 1130
rect 2320 773 2322 1007
rect 2368 773 2370 1007
rect 2320 720 2370 773
rect 2490 1032 2540 1060
rect 2490 798 2492 1032
rect 2538 798 2540 1032
rect 2490 670 2540 798
rect 2660 1007 2710 1130
rect 2660 773 2662 1007
rect 2708 773 2710 1007
rect 2830 1032 2880 1060
rect 2830 798 2832 1032
rect 2878 798 2880 1032
rect 2830 780 2880 798
rect 3000 1007 3050 1130
rect 2660 720 2710 773
rect 2810 776 2910 780
rect 2810 724 2834 776
rect 2886 724 2910 776
rect 2810 720 2910 724
rect 3000 773 3002 1007
rect 3048 773 3050 1007
rect 3000 720 3050 773
rect 2830 670 2880 720
rect 110 663 400 670
rect 110 617 327 663
rect 373 617 400 663
rect 110 610 400 617
rect 450 610 2880 670
rect 110 318 160 610
rect 210 516 310 520
rect 210 464 234 516
rect 286 464 310 516
rect 210 460 310 464
rect 450 490 500 610
rect 790 490 840 610
rect 1130 490 1180 610
rect 1470 490 1520 610
rect 1810 490 1860 610
rect 2150 490 2200 610
rect 2490 490 2540 610
rect 2830 490 2880 610
rect 450 430 2880 490
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 450 318 500 430
rect 450 272 452 318
rect 498 272 500 318
rect 450 210 500 272
rect 620 318 670 380
rect 620 272 622 318
rect 668 272 670 318
rect 620 140 670 272
rect 790 318 840 430
rect 790 272 792 318
rect 838 272 840 318
rect 790 210 840 272
rect 960 318 1010 380
rect 960 272 962 318
rect 1008 272 1010 318
rect 960 140 1010 272
rect 1130 318 1180 430
rect 1130 272 1132 318
rect 1178 272 1180 318
rect 1130 210 1180 272
rect 1300 318 1350 380
rect 1300 272 1302 318
rect 1348 272 1350 318
rect 1300 140 1350 272
rect 1470 318 1520 430
rect 1470 272 1472 318
rect 1518 272 1520 318
rect 1470 210 1520 272
rect 1640 318 1690 380
rect 1640 272 1642 318
rect 1688 272 1690 318
rect 1640 140 1690 272
rect 1810 318 1860 430
rect 1810 272 1812 318
rect 1858 272 1860 318
rect 1810 210 1860 272
rect 1980 318 2030 380
rect 1980 272 1982 318
rect 2028 272 2030 318
rect 1980 140 2030 272
rect 2150 318 2200 430
rect 2150 272 2152 318
rect 2198 272 2200 318
rect 2150 210 2200 272
rect 2320 318 2370 380
rect 2320 272 2322 318
rect 2368 272 2370 318
rect 2320 140 2370 272
rect 2490 318 2540 430
rect 2490 272 2492 318
rect 2538 272 2540 318
rect 2490 210 2540 272
rect 2660 318 2710 380
rect 2660 272 2662 318
rect 2708 272 2710 318
rect 2660 140 2710 272
rect 2830 318 2880 430
rect 2830 272 2832 318
rect 2878 272 2880 318
rect 2830 210 2880 272
rect 3000 318 3050 380
rect 3000 272 3002 318
rect 3048 272 3050 318
rect 3000 140 3050 272
rect 0 118 3160 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1312 118
rect 1358 72 1552 118
rect 1598 72 1792 118
rect 1838 72 2032 118
rect 2078 72 2272 118
rect 2318 72 2512 118
rect 2558 72 2752 118
rect 2798 72 3160 118
rect 0 0 3160 72
<< via1 >>
rect 2834 724 2886 776
rect 234 513 286 516
rect 234 467 237 513
rect 237 467 283 513
rect 283 467 286 513
rect 234 464 286 467
<< metal2 >>
rect 2810 776 2910 790
rect 2810 724 2834 776
rect 2886 724 2910 776
rect 2810 710 2910 724
rect 220 520 300 530
rect 210 516 310 520
rect 210 464 234 516
rect 286 464 310 516
rect 210 460 310 464
rect 220 450 300 460
<< labels >>
rlabel via1 s 234 464 286 516 4 A
port 1 nsew signal input
rlabel via1 s 2834 724 2886 776 4 Y
port 2 nsew signal output
rlabel metal1 s 280 720 330 1270 4 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 620 720 670 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 960 720 1010 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1300 720 1350 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1640 720 1690 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1980 720 2030 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2320 720 2370 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2660 720 2710 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3000 720 3050 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 1130 3160 1270 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 620 0 670 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 960 0 1010 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1300 0 1350 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1640 0 1690 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1980 0 2030 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2320 0 2370 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2660 0 2710 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3000 0 3050 380 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 0 3160 140 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal2 s 220 450 300 530 1 A
port 1 nsew signal input
rlabel metal2 s 210 460 310 520 1 A
port 1 nsew signal input
rlabel metal1 s 210 460 310 520 1 A
port 1 nsew signal input
rlabel metal2 s 2810 710 2910 790 1 Y
port 2 nsew signal output
rlabel metal1 s 450 210 500 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 790 210 840 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 1130 210 1180 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 1470 210 1520 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 1810 210 1860 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 2150 210 2200 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 2490 210 2540 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 450 430 2880 490 1 Y
port 2 nsew signal output
rlabel metal1 s 450 610 2880 670 1 Y
port 2 nsew signal output
rlabel metal1 s 2830 210 2880 1060 1 Y
port 2 nsew signal output
rlabel metal1 s 2810 720 2910 780 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3160 1270
string GDS_END 95644
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 78844
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
