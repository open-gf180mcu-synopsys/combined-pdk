VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__asig_5p0
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_fd_io__asig_5p0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN ASIG5V
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1200.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.340 134.370 17.880 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 51.440 134.370 53.980 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 57.120 134.370 59.660 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 21.020 134.370 23.560 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 45.760 134.370 48.300 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 40.080 134.370 42.620 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 32.380 134.370 34.920 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 26.700 134.370 29.240 350.000 ;
    END
  END ASIG5V
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 70.820 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.820 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 4.180 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 5.570 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 5.570 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 5.570 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 5.570 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 4.180 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 4.180 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 4.180 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 4.180 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 4.180 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 4.180 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 4.180 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 73.660 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 73.660 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 1.340 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 1.340 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 1.340 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 1.340 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.340 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.340 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 1.340 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.340 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.340 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.340 117.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 4.930 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 4.930 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 4.030 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 4.030 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 134.070 15.040 348.390 ;
        RECT 18.180 134.070 20.720 348.390 ;
        RECT 23.860 134.070 26.400 348.390 ;
        RECT 29.540 134.070 32.080 348.390 ;
        RECT 35.220 134.070 39.780 348.390 ;
        RECT 42.920 134.070 45.460 348.390 ;
        RECT 48.600 134.070 51.140 348.390 ;
        RECT 54.280 134.070 56.820 348.390 ;
        RECT 59.960 134.070 75.000 348.390 ;
        RECT 0.000 0.000 75.000 134.070 ;
      LAYER Metal3 ;
        RECT 3.140 342.800 71.860 348.390 ;
        RECT 5.980 332.200 69.020 342.800 ;
        RECT 3.140 324.200 71.860 332.200 ;
        RECT 2.800 318.800 72.200 324.200 ;
        RECT 3.140 302.800 71.860 308.200 ;
        RECT 7.370 292.200 69.020 302.800 ;
        RECT 3.140 286.800 71.860 292.200 ;
        RECT 7.370 262.800 69.020 286.800 ;
        RECT 2.800 246.800 72.200 252.200 ;
        RECT 3.140 230.800 71.860 246.800 ;
        RECT 5.980 204.200 69.020 230.800 ;
        RECT 3.140 198.800 71.860 204.200 ;
        RECT 5.980 132.200 69.020 198.800 ;
        RECT 3.140 126.800 71.860 132.200 ;
        RECT 5.980 116.200 69.020 126.800 ;
        RECT 3.140 68.200 71.860 116.200 ;
        RECT 1.000 0.000 74.000 68.200 ;
  END
END gf180mcu_fd_io__asig_5p0
END LIBRARY

