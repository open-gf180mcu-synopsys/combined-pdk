magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
use pmos_5p043105899832106_64x8m81  pmos_5p043105899832106_64x8m81_0
timestamp 1750858719
transform 1 0 -31 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 405564
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 405058
<< end >>
