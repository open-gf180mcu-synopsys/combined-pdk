magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 352 534 870
<< pwell >>
rect -86 -86 534 352
<< metal1 >>
rect 0 724 448 844
rect 50 472 96 724
rect 244 461 316 678
rect 50 60 96 232
rect 0 -60 448 60
<< obsm1 >>
rect 175 267 320 314
rect 274 106 320 267
<< labels >>
rlabel metal1 s 244 461 316 678 6 Z
port 1 nsew default output
rlabel metal1 s 50 472 96 724 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 724 448 844 6 VDD
port 2 nsew power bidirectional abutment
rlabel nwell s -86 352 534 870 6 VNW
port 3 nsew power bidirectional
rlabel pwell s -86 -86 534 352 6 VPW
port 4 nsew ground bidirectional
rlabel metal1 s 0 -60 448 60 8 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 50 60 96 232 6 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string LEFclass core TIEHIGH
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 318162
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 316076
<< end >>
