magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 730 1660
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 470 210 530 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 470 1110 530 1450
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 470 380
rect 530 318 630 380
rect 530 272 562 318
rect 608 272 630 318
rect 530 210 630 272
<< pdiff >>
rect 90 1397 190 1450
rect 90 1163 112 1397
rect 158 1163 190 1397
rect 90 1110 190 1163
rect 250 1397 360 1450
rect 250 1163 282 1397
rect 328 1163 360 1397
rect 250 1110 360 1163
rect 420 1110 470 1450
rect 530 1397 630 1450
rect 530 1163 562 1397
rect 608 1163 630 1397
rect 530 1110 630 1163
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 562 272 608 318
<< pdiffc >>
rect 112 1163 158 1397
rect 282 1163 328 1397
rect 562 1163 608 1397
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 470 1450 530 1500
rect 190 540 250 1110
rect 360 1060 420 1110
rect 300 1038 420 1060
rect 300 992 322 1038
rect 368 992 420 1038
rect 300 970 420 992
rect 470 1060 530 1110
rect 470 1038 630 1060
rect 470 992 562 1038
rect 608 992 630 1038
rect 470 970 630 992
rect 190 518 310 540
rect 190 472 232 518
rect 278 472 310 518
rect 190 450 310 472
rect 190 380 250 450
rect 360 380 420 970
rect 470 508 630 530
rect 470 462 562 508
rect 608 462 630 508
rect 470 440 630 462
rect 470 380 530 440
rect 190 160 250 210
rect 360 160 420 210
rect 470 160 530 210
<< polycontact >>
rect 322 992 368 1038
rect 562 992 608 1038
rect 232 472 278 518
rect 562 462 608 508
<< metal1 >>
rect 0 1588 730 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 730 1588
rect 0 1520 730 1542
rect 110 1397 160 1450
rect 110 1163 112 1397
rect 158 1163 160 1397
rect 110 1160 160 1163
rect 100 1110 160 1160
rect 280 1397 330 1520
rect 280 1163 282 1397
rect 328 1163 330 1397
rect 280 1110 330 1163
rect 560 1397 610 1450
rect 560 1163 562 1397
rect 608 1163 610 1397
rect 560 1160 610 1163
rect 440 1110 610 1160
rect 100 910 150 1110
rect 290 1038 390 1040
rect 290 1036 322 1038
rect 290 984 314 1036
rect 368 992 390 1038
rect 366 984 390 992
rect 290 980 390 984
rect 70 906 170 910
rect 70 854 94 906
rect 146 854 170 906
rect 70 850 170 854
rect 100 430 150 850
rect 440 780 490 1110
rect 540 1038 640 1040
rect 540 992 562 1038
rect 608 1036 640 1038
rect 540 984 564 992
rect 616 984 640 1036
rect 540 980 640 984
rect 410 776 520 780
rect 410 724 434 776
rect 486 724 520 776
rect 410 720 520 724
rect 200 518 300 520
rect 200 516 232 518
rect 200 464 224 516
rect 278 472 300 518
rect 276 464 300 472
rect 200 460 300 464
rect 100 380 160 430
rect 440 380 490 720
rect 540 516 640 520
rect 540 508 564 516
rect 540 462 562 508
rect 616 464 640 516
rect 608 462 640 464
rect 540 460 640 462
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 440 330 610 380
rect 280 272 282 318
rect 328 272 330 318
rect 280 140 330 272
rect 560 318 610 330
rect 560 272 562 318
rect 608 272 610 318
rect 560 210 610 272
rect 0 118 730 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 730 118
rect 0 0 730 72
<< via1 >>
rect 314 992 322 1036
rect 322 992 366 1036
rect 314 984 366 992
rect 94 854 146 906
rect 564 992 608 1036
rect 608 992 616 1036
rect 564 984 616 992
rect 434 724 486 776
rect 224 472 232 516
rect 232 472 276 516
rect 224 464 276 472
rect 564 508 616 516
rect 564 464 608 508
rect 608 464 616 508
<< metal2 >>
rect 290 1036 390 1050
rect 290 984 314 1036
rect 366 984 390 1036
rect 290 970 390 984
rect 540 1036 640 1050
rect 540 984 564 1036
rect 616 984 640 1036
rect 540 970 640 984
rect 70 910 170 920
rect 560 910 620 970
rect 70 906 620 910
rect 70 854 94 906
rect 146 854 620 906
rect 70 850 620 854
rect 70 840 170 850
rect 410 776 510 790
rect 410 724 434 776
rect 486 724 510 776
rect 410 710 510 724
rect 200 520 300 530
rect 540 520 640 530
rect 200 516 640 520
rect 200 464 224 516
rect 276 464 564 516
rect 616 464 640 516
rect 200 460 640 464
rect 200 450 300 460
rect 540 450 640 460
<< labels >>
rlabel via1 s 314 984 366 1036 4 A
port 1 nsew signal input
rlabel via1 s 434 724 486 776 4 Y
port 2 nsew signal output
rlabel via1 s 564 464 616 516 4 EN
port 3 nsew signal input
rlabel metal1 s 280 1110 330 1660 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 1520 730 1660 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 0 730 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal2 s 290 970 390 1050 1 A
port 1 nsew signal input
rlabel metal1 s 290 980 390 1040 1 A
port 1 nsew signal input
rlabel via1 s 224 464 276 516 1 EN
port 3 nsew signal input
rlabel metal2 s 200 450 300 530 1 EN
port 3 nsew signal input
rlabel metal2 s 200 460 640 520 1 EN
port 3 nsew signal input
rlabel metal2 s 540 450 640 530 1 EN
port 3 nsew signal input
rlabel metal1 s 200 460 300 520 1 EN
port 3 nsew signal input
rlabel metal1 s 540 460 640 520 1 EN
port 3 nsew signal input
rlabel metal2 s 410 710 510 790 1 Y
port 2 nsew signal output
rlabel metal1 s 440 330 490 1160 1 Y
port 2 nsew signal output
rlabel metal1 s 410 720 520 780 1 Y
port 2 nsew signal output
rlabel metal1 s 440 1110 610 1160 1 Y
port 2 nsew signal output
rlabel metal1 s 560 210 610 380 1 Y
port 2 nsew signal output
rlabel metal1 s 440 330 610 380 1 Y
port 2 nsew signal output
rlabel metal1 s 560 1110 610 1450 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 730 1660
string GDS_END 515706
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 509812
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
