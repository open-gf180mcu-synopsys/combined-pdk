magic
tech gf180mcuA
magscale 1 5
timestamp 1750858719
<< metal1 >>
rect 0 565 220 635
rect 55 360 80 565
rect 140 195 165 200
rect 130 193 180 195
rect 55 70 80 190
rect 130 167 142 193
rect 168 167 180 193
rect 130 165 180 167
rect 140 105 165 165
rect 0 0 220 70
<< via1 >>
rect 142 167 168 193
<< obsm1 >>
rect 140 325 165 530
rect 115 300 165 325
<< metal2 >>
rect 130 193 180 200
rect 130 167 142 193
rect 168 167 180 193
rect 130 160 180 167
<< labels >>
rlabel metal1 s 55 360 80 635 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 565 220 635 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 55 0 80 190 6 VSS
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 0 220 70 6 VSS
port 3 nsew ground bidirectional abutment
rlabel via1 s 142 167 168 193 6 Y
port 1 nsew signal output
rlabel metal2 s 130 160 180 200 6 Y
port 1 nsew signal output
rlabel metal1 s 140 105 165 200 6 Y
port 1 nsew signal output
rlabel metal1 s 130 165 180 195 6 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 220 635
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 372648
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 370094
<< end >>
