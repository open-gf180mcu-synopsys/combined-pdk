magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect -86 377 2774 870
rect -86 352 2158 377
rect 2378 352 2774 377
<< pwell >>
rect 2158 352 2378 377
rect -86 -86 2774 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 608 93 728 165
rect 832 93 952 165
rect 1016 93 1136 165
rect 1384 93 1504 165
rect 1568 93 1688 165
rect 1828 68 1948 232
rect 2052 68 2172 232
rect 2364 68 2484 232
<< mvpmos >>
rect 144 567 244 639
rect 358 567 458 639
rect 618 527 718 639
rect 832 527 932 639
rect 1036 527 1136 639
rect 1384 527 1484 639
rect 1588 527 1688 639
rect 1848 497 1948 716
rect 2072 497 2172 716
rect 2364 497 2464 716
<< mvndiff >>
rect 2232 244 2304 257
rect 2232 232 2245 244
rect 1748 165 1828 232
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 608 165
rect 468 106 497 152
rect 543 106 608 152
rect 468 93 608 106
rect 728 152 832 165
rect 728 106 757 152
rect 803 106 832 152
rect 728 93 832 106
rect 952 93 1016 165
rect 1136 152 1224 165
rect 1136 106 1165 152
rect 1211 106 1224 152
rect 1136 93 1224 106
rect 1296 152 1384 165
rect 1296 106 1309 152
rect 1355 106 1384 152
rect 1296 93 1384 106
rect 1504 93 1568 165
rect 1688 152 1828 165
rect 1688 106 1717 152
rect 1763 106 1828 152
rect 1688 93 1828 106
rect 1748 68 1828 93
rect 1948 152 2052 232
rect 1948 106 1977 152
rect 2023 106 2052 152
rect 1948 68 2052 106
rect 2172 198 2245 232
rect 2291 232 2304 244
rect 2291 198 2364 232
rect 2172 68 2364 198
rect 2484 152 2572 232
rect 2484 106 2513 152
rect 2559 106 2572 152
rect 2484 68 2572 106
<< mvpdiff >>
rect 1750 703 1848 716
rect 1750 639 1763 703
rect 56 626 144 639
rect 56 580 69 626
rect 115 580 144 626
rect 56 567 144 580
rect 244 567 358 639
rect 458 626 618 639
rect 458 580 487 626
rect 533 580 618 626
rect 458 567 618 580
rect 538 527 618 567
rect 718 626 832 639
rect 718 580 757 626
rect 803 580 832 626
rect 718 527 832 580
rect 932 586 1036 639
rect 932 540 961 586
rect 1007 540 1036 586
rect 932 527 1036 540
rect 1136 626 1224 639
rect 1136 580 1165 626
rect 1211 580 1224 626
rect 1136 527 1224 580
rect 1296 626 1384 639
rect 1296 580 1309 626
rect 1355 580 1384 626
rect 1296 527 1384 580
rect 1484 586 1588 639
rect 1484 540 1513 586
rect 1559 540 1588 586
rect 1484 527 1588 540
rect 1688 563 1763 639
rect 1809 563 1848 703
rect 1688 527 1848 563
rect 1758 497 1848 527
rect 1948 639 2072 716
rect 1948 593 1997 639
rect 2043 593 2072 639
rect 1948 497 2072 593
rect 2172 497 2364 716
rect 2464 689 2552 716
rect 2464 643 2493 689
rect 2539 643 2552 689
rect 2464 497 2552 643
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 497 106 543 152
rect 757 106 803 152
rect 1165 106 1211 152
rect 1309 106 1355 152
rect 1717 106 1763 152
rect 1977 106 2023 152
rect 2245 198 2291 244
rect 2513 106 2559 152
<< mvpdiffc >>
rect 69 580 115 626
rect 487 580 533 626
rect 757 580 803 626
rect 961 540 1007 586
rect 1165 580 1211 626
rect 1309 580 1355 626
rect 1513 540 1559 586
rect 1763 563 1809 703
rect 1997 593 2043 639
rect 2493 643 2539 689
<< polysilicon >>
rect 1848 716 1948 760
rect 2072 716 2172 760
rect 2364 716 2464 760
rect 144 639 244 683
rect 358 639 458 683
rect 618 639 718 683
rect 832 639 932 683
rect 1036 639 1136 683
rect 1384 639 1484 683
rect 1588 639 1688 683
rect 144 526 244 567
rect 144 480 185 526
rect 231 480 244 526
rect 144 209 244 480
rect 358 375 458 567
rect 358 329 386 375
rect 432 329 458 375
rect 358 209 458 329
rect 618 244 718 527
rect 618 209 640 244
rect 124 165 244 209
rect 348 165 468 209
rect 608 198 640 209
rect 686 209 718 244
rect 832 338 932 527
rect 832 292 857 338
rect 903 292 932 338
rect 832 209 932 292
rect 1036 390 1136 527
rect 1036 344 1058 390
rect 1104 344 1136 390
rect 1036 209 1136 344
rect 686 198 728 209
rect 608 165 728 198
rect 832 165 952 209
rect 1016 165 1136 209
rect 1384 465 1484 527
rect 1384 325 1406 465
rect 1452 325 1484 465
rect 1384 209 1484 325
rect 1588 415 1688 527
rect 1588 369 1629 415
rect 1675 369 1688 415
rect 1588 209 1688 369
rect 1848 348 1948 497
rect 1828 313 1948 348
rect 1828 267 1851 313
rect 1897 267 1948 313
rect 2072 416 2172 497
rect 2072 370 2093 416
rect 2139 370 2172 416
rect 2072 288 2172 370
rect 1828 232 1948 267
rect 2052 232 2172 288
rect 2364 419 2464 497
rect 2364 373 2377 419
rect 2423 373 2464 419
rect 2364 288 2464 373
rect 1384 165 1504 209
rect 1568 165 1688 209
rect 124 49 244 93
rect 348 49 468 93
rect 608 49 728 93
rect 832 49 952 93
rect 1016 49 1136 93
rect 1384 49 1504 93
rect 1568 49 1688 93
rect 2364 232 2484 288
rect 1828 24 1948 68
rect 2052 24 2172 68
rect 2364 24 2484 68
<< polycontact >>
rect 185 480 231 526
rect 386 329 432 375
rect 640 198 686 244
rect 857 292 903 338
rect 1058 344 1104 390
rect 1406 325 1452 465
rect 1629 369 1675 415
rect 1851 267 1897 313
rect 2093 370 2139 416
rect 2377 373 2423 419
<< metal1 >>
rect 0 724 2688 844
rect 69 626 115 639
rect 474 626 546 724
rect 474 580 487 626
rect 533 580 546 626
rect 744 632 1224 678
rect 744 626 816 632
rect 744 580 757 626
rect 803 580 816 626
rect 1152 626 1224 632
rect 69 244 115 580
rect 948 540 961 586
rect 1007 540 1020 586
rect 1152 580 1165 626
rect 1211 580 1224 626
rect 1309 626 1355 724
rect 1752 703 1820 724
rect 1309 568 1355 580
rect 1406 632 1700 678
rect 174 526 872 531
rect 174 480 185 526
rect 231 480 872 526
rect 174 477 872 480
rect 826 430 872 477
rect 948 522 1020 540
rect 1406 522 1452 632
rect 948 476 1452 522
rect 354 375 780 419
rect 826 390 1124 430
rect 826 384 1058 390
rect 354 329 386 375
rect 432 365 780 375
rect 432 329 445 365
rect 354 291 445 329
rect 734 338 780 365
rect 1035 344 1058 384
rect 1104 344 1124 390
rect 734 292 857 338
rect 903 292 954 338
rect 1035 319 1124 344
rect 734 291 954 292
rect 1176 245 1222 476
rect 1406 465 1452 476
rect 1406 307 1452 325
rect 1502 540 1513 586
rect 1559 540 1570 586
rect 1502 245 1570 540
rect 1654 513 1700 632
rect 1752 563 1763 703
rect 1809 563 1820 703
rect 2493 689 2539 724
rect 1914 639 2443 648
rect 1914 593 1997 639
rect 2043 593 2443 639
rect 2493 603 2539 643
rect 1914 584 2443 593
rect 2376 536 2443 584
rect 1654 466 2290 513
rect 2376 472 2552 536
rect 2244 419 2290 466
rect 1617 416 2153 419
rect 1617 415 2093 416
rect 1617 369 1629 415
rect 1675 370 2093 415
rect 2139 370 2153 416
rect 2244 373 2377 419
rect 2423 373 2434 419
rect 2244 372 2434 373
rect 1675 369 2153 370
rect 1617 365 2153 369
rect 2488 316 2552 472
rect 1840 267 1851 313
rect 1897 267 1908 313
rect 1840 245 1908 267
rect 69 198 640 244
rect 686 198 699 244
rect 746 198 1222 245
rect 1298 198 1908 245
rect 2234 244 2552 316
rect 2234 198 2245 244
rect 2291 198 2552 244
rect 261 152 330 198
rect 746 152 814 198
rect 1298 152 1366 198
rect 38 106 49 152
rect 95 106 106 152
rect 261 106 273 152
rect 319 106 330 152
rect 486 106 497 152
rect 543 106 554 152
rect 746 106 757 152
rect 803 106 814 152
rect 1154 106 1165 152
rect 1211 106 1222 152
rect 1298 106 1309 152
rect 1355 106 1366 152
rect 1706 106 1717 152
rect 1763 106 1774 152
rect 1948 106 1977 152
rect 2023 106 2513 152
rect 2559 106 2572 152
rect 38 60 106 106
rect 486 60 554 106
rect 1154 60 1222 106
rect 1706 60 1774 106
rect 0 -60 2688 60
<< labels >>
flabel metal1 s 1617 365 2153 419 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 2688 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1706 60 1774 152 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 1914 584 2443 648 0 FreeSans 400 0 0 0 ZN
port 4 nsew default output
flabel metal1 s 354 365 780 419 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 174 477 872 531 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 734 338 780 365 1 A1
port 1 nsew default input
rlabel metal1 s 354 338 445 365 1 A1
port 1 nsew default input
rlabel metal1 s 734 291 954 338 1 A1
port 1 nsew default input
rlabel metal1 s 354 291 445 338 1 A1
port 1 nsew default input
rlabel metal1 s 826 430 872 477 1 A2
port 2 nsew default input
rlabel metal1 s 826 384 1124 430 1 A2
port 2 nsew default input
rlabel metal1 s 1035 319 1124 384 1 A2
port 2 nsew default input
rlabel metal1 s 2376 536 2443 584 1 ZN
port 4 nsew default output
rlabel metal1 s 2376 472 2552 536 1 ZN
port 4 nsew default output
rlabel metal1 s 2488 316 2552 472 1 ZN
port 4 nsew default output
rlabel metal1 s 2234 198 2552 316 1 ZN
port 4 nsew default output
rlabel metal1 s 2493 603 2539 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1752 603 1820 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1309 603 1355 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 474 603 546 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1752 580 1820 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1309 580 1355 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 474 580 546 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1752 568 1820 580 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1309 568 1355 580 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1752 563 1820 568 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1154 60 1222 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2688 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2688 784
string GDS_END 341068
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 334956
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
