magic
tech gf180mcuA
timestamp 1750858719
<< properties >>
string GDS_END 375394
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 371486
<< end >>
