magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 630 1280 1270
<< nmos >>
rect 190 210 250 380
rect 360 210 420 380
rect 490 210 550 380
rect 720 210 780 380
rect 850 210 910 380
rect 1020 210 1080 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 490 720 550 1060
rect 720 720 780 1060
rect 850 720 910 1060
rect 1020 720 1080 1060
<< ndiff >>
rect 580 380 680 390
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 360 380
rect 250 272 282 318
rect 328 272 360 318
rect 250 210 360 272
rect 420 210 490 380
rect 550 370 720 380
rect 550 230 612 370
rect 658 230 720 370
rect 550 210 720 230
rect 780 210 850 380
rect 910 318 1020 380
rect 910 272 942 318
rect 988 272 1020 318
rect 910 210 1020 272
rect 1080 318 1180 380
rect 1080 272 1112 318
rect 1158 272 1180 318
rect 1080 210 1180 272
<< pdiff >>
rect 90 1023 190 1060
rect 90 977 112 1023
rect 158 977 190 1023
rect 90 720 190 977
rect 250 1023 360 1060
rect 250 977 282 1023
rect 328 977 360 1023
rect 250 720 360 977
rect 420 720 490 1060
rect 550 1023 720 1060
rect 550 977 612 1023
rect 658 977 720 1023
rect 550 720 720 977
rect 780 720 850 1060
rect 910 1023 1020 1060
rect 910 977 942 1023
rect 988 977 1020 1023
rect 910 720 1020 977
rect 1080 1023 1180 1060
rect 1080 977 1112 1023
rect 1158 977 1180 1023
rect 1080 720 1180 977
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 612 230 658 370
rect 942 272 988 318
rect 1112 272 1158 318
<< pdiffc >>
rect 112 977 158 1023
rect 282 977 328 1023
rect 612 977 658 1023
rect 942 977 988 1023
rect 1112 977 1158 1023
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 300 118 450 140
rect 300 72 352 118
rect 398 72 450 118
rect 300 50 450 72
rect 540 118 690 140
rect 540 72 592 118
rect 638 72 690 118
rect 540 50 690 72
rect 780 118 930 140
rect 780 72 832 118
rect 878 72 930 118
rect 780 50 930 72
rect 1020 118 1170 140
rect 1020 72 1072 118
rect 1118 72 1170 118
rect 1020 50 1170 72
<< nsubdiff >>
rect 60 1198 210 1220
rect 60 1152 112 1198
rect 158 1152 210 1198
rect 60 1130 210 1152
rect 300 1198 450 1220
rect 300 1152 352 1198
rect 398 1152 450 1198
rect 300 1130 450 1152
rect 540 1198 690 1220
rect 540 1152 592 1198
rect 638 1152 690 1198
rect 540 1130 690 1152
rect 780 1198 930 1220
rect 780 1152 832 1198
rect 878 1152 930 1198
rect 780 1130 930 1152
rect 1020 1198 1170 1220
rect 1020 1152 1072 1198
rect 1118 1152 1170 1198
rect 1020 1130 1170 1152
<< psubdiffcont >>
rect 112 72 158 118
rect 352 72 398 118
rect 592 72 638 118
rect 832 72 878 118
rect 1072 72 1118 118
<< nsubdiffcont >>
rect 112 1152 158 1198
rect 352 1152 398 1198
rect 592 1152 638 1198
rect 832 1152 878 1198
rect 1072 1152 1118 1198
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 490 1060 550 1110
rect 720 1060 780 1110
rect 850 1060 910 1110
rect 1020 1060 1080 1110
rect 190 540 250 720
rect 360 700 420 720
rect 310 673 420 700
rect 310 627 337 673
rect 383 627 420 673
rect 310 600 420 627
rect 490 700 550 720
rect 720 700 780 720
rect 850 700 910 720
rect 1020 700 1080 720
rect 490 673 630 700
rect 490 627 557 673
rect 603 627 630 673
rect 490 600 630 627
rect 700 673 800 700
rect 700 627 727 673
rect 773 627 800 673
rect 850 650 1080 700
rect 700 600 800 627
rect 190 513 350 540
rect 190 467 277 513
rect 323 510 350 513
rect 323 467 420 510
rect 190 440 420 467
rect 190 380 250 440
rect 360 380 420 440
rect 490 380 550 600
rect 1020 540 1080 650
rect 600 520 700 540
rect 600 513 780 520
rect 600 467 627 513
rect 673 467 780 513
rect 910 513 1080 540
rect 910 490 937 513
rect 600 440 780 467
rect 720 380 780 440
rect 850 467 937 490
rect 983 467 1080 513
rect 850 440 1080 467
rect 850 380 910 440
rect 1020 380 1080 440
rect 190 160 250 210
rect 360 160 420 210
rect 490 160 550 210
rect 720 160 780 210
rect 850 160 910 210
rect 1020 160 1080 210
<< polycontact >>
rect 337 627 383 673
rect 557 627 603 673
rect 727 627 773 673
rect 277 467 323 513
rect 627 467 673 513
rect 937 467 983 513
<< metal1 >>
rect 0 1198 1280 1270
rect 0 1152 112 1198
rect 158 1152 352 1198
rect 398 1152 592 1198
rect 638 1152 832 1198
rect 878 1152 1072 1198
rect 1118 1152 1280 1198
rect 0 1130 1280 1152
rect 110 1023 160 1060
rect 110 977 112 1023
rect 158 977 160 1023
rect 110 680 160 977
rect 280 1023 330 1130
rect 280 977 282 1023
rect 328 977 330 1023
rect 280 940 330 977
rect 610 1023 660 1060
rect 610 977 612 1023
rect 658 977 660 1023
rect 610 970 660 977
rect 600 906 660 970
rect 940 1023 990 1130
rect 940 977 942 1023
rect 988 977 990 1023
rect 940 940 990 977
rect 1110 1023 1160 1060
rect 1110 977 1112 1023
rect 1158 977 1160 1023
rect 600 854 604 906
rect 656 854 660 906
rect 600 830 660 854
rect 1110 780 1160 977
rect 550 730 1160 780
rect 110 673 480 680
rect 110 627 337 673
rect 383 627 480 673
rect 110 620 480 627
rect 110 318 160 620
rect 420 520 480 620
rect 550 673 610 730
rect 550 627 557 673
rect 603 627 610 673
rect 550 600 610 627
rect 700 676 800 680
rect 700 624 724 676
rect 776 624 800 676
rect 700 620 800 624
rect 250 516 350 520
rect 250 464 274 516
rect 326 464 350 516
rect 250 460 350 464
rect 420 513 700 520
rect 420 467 627 513
rect 673 467 700 513
rect 420 460 700 467
rect 910 516 1010 520
rect 910 464 934 516
rect 986 464 1010 516
rect 910 460 1010 464
rect 600 386 660 410
rect 110 272 112 318
rect 158 272 160 318
rect 110 210 160 272
rect 280 318 330 380
rect 280 272 282 318
rect 328 272 330 318
rect 600 334 604 386
rect 656 370 660 386
rect 600 300 612 334
rect 280 140 330 272
rect 610 230 612 300
rect 658 230 660 370
rect 610 210 660 230
rect 940 318 990 380
rect 940 272 942 318
rect 988 272 990 318
rect 940 140 990 272
rect 1110 318 1160 730
rect 1110 272 1112 318
rect 1158 272 1160 318
rect 1110 210 1160 272
rect 0 118 1280 140
rect 0 72 112 118
rect 158 72 352 118
rect 398 72 592 118
rect 638 72 832 118
rect 878 72 1072 118
rect 1118 72 1280 118
rect 0 0 1280 72
<< via1 >>
rect 604 854 656 906
rect 724 673 776 676
rect 724 627 727 673
rect 727 627 773 673
rect 773 627 776 673
rect 724 624 776 627
rect 274 513 326 516
rect 274 467 277 513
rect 277 467 323 513
rect 323 467 326 513
rect 274 464 326 467
rect 934 513 986 516
rect 934 467 937 513
rect 937 467 983 513
rect 983 467 986 513
rect 934 464 986 467
rect 604 370 656 386
rect 604 334 612 370
rect 612 334 656 370
<< metal2 >>
rect 600 920 660 970
rect 590 906 670 920
rect 590 854 604 906
rect 656 854 670 906
rect 590 840 670 854
rect 590 830 660 840
rect 270 530 330 540
rect 260 516 340 530
rect 260 464 274 516
rect 326 464 340 516
rect 260 450 340 464
rect 270 260 330 450
rect 590 400 650 830
rect 720 690 790 700
rect 710 676 800 690
rect 710 624 724 676
rect 776 624 800 676
rect 710 610 800 624
rect 720 600 800 610
rect 580 386 680 400
rect 580 334 604 386
rect 656 334 680 386
rect 580 320 680 334
rect 740 260 800 600
rect 930 530 990 540
rect 920 520 1000 530
rect 910 516 1010 520
rect 910 464 934 516
rect 986 464 1010 516
rect 910 460 1010 464
rect 920 450 1000 460
rect 930 440 990 450
rect 270 200 800 260
<< labels >>
rlabel via1 s 724 624 776 676 4 A
port 1 nsew signal input
rlabel via1 s 934 464 986 516 4 B
port 2 nsew signal input
rlabel via1 s 604 334 656 386 4 Y
port 3 nsew signal output
rlabel metal1 s 280 940 330 1270 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 280 0 330 380 4 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 940 940 990 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 1130 1280 1270 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 940 0 990 380 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1280 140 1 VSS
port 5 nsew ground bidirectional abutment
rlabel via1 s 274 464 326 516 1 A
port 1 nsew signal input
rlabel metal2 s 270 200 330 540 1 A
port 1 nsew signal input
rlabel metal2 s 260 450 340 530 1 A
port 1 nsew signal input
rlabel metal2 s 270 200 800 260 1 A
port 1 nsew signal input
rlabel metal2 s 720 600 790 700 1 A
port 1 nsew signal input
rlabel metal2 s 740 200 800 690 1 A
port 1 nsew signal input
rlabel metal2 s 710 610 800 690 1 A
port 1 nsew signal input
rlabel metal1 s 250 460 350 520 1 A
port 1 nsew signal input
rlabel metal1 s 700 620 800 680 1 A
port 1 nsew signal input
rlabel metal2 s 930 440 990 540 1 B
port 2 nsew signal input
rlabel metal2 s 920 450 1000 530 1 B
port 2 nsew signal input
rlabel metal2 s 910 460 1010 520 1 B
port 2 nsew signal input
rlabel metal1 s 910 460 1010 520 1 B
port 2 nsew signal input
rlabel via1 s 604 854 656 906 1 Y
port 3 nsew signal output
rlabel metal2 s 590 320 650 920 1 Y
port 3 nsew signal output
rlabel metal2 s 600 830 660 970 1 Y
port 3 nsew signal output
rlabel metal2 s 590 840 670 920 1 Y
port 3 nsew signal output
rlabel metal2 s 580 320 680 400 1 Y
port 3 nsew signal output
rlabel metal1 s 600 830 660 970 1 Y
port 3 nsew signal output
rlabel metal1 s 610 830 660 1060 1 Y
port 3 nsew signal output
rlabel metal1 s 610 210 660 410 1 Y
port 3 nsew signal output
rlabel metal1 s 600 300 660 410 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1280 1270
string GDS_END 387188
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp9t3v3/gds/gf180mcu_osu_sc_gp9t3v3.gds
string GDS_START 378990
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp9t3v3
string LEFsymmetry X Y
<< end >>
