magic
tech gf180mcuA
magscale 1 10
timestamp 1750858719
<< nwell >>
rect 0 1020 1070 1660
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
rect 500 210 560 380
rect 610 210 670 380
<< pmos >>
rect 190 1110 250 1450
rect 360 1110 420 1450
rect 530 1110 590 1450
rect 700 1110 760 1450
<< ndiff >>
rect 120 318 220 380
rect 120 272 142 318
rect 188 272 220 318
rect 120 210 220 272
rect 280 210 330 380
rect 390 318 500 380
rect 390 272 422 318
rect 468 272 500 318
rect 390 210 500 272
rect 560 210 610 380
rect 670 318 770 380
rect 670 272 702 318
rect 748 272 770 318
rect 670 210 770 272
<< pdiff >>
rect 90 1425 190 1450
rect 90 1285 112 1425
rect 158 1285 190 1425
rect 90 1110 190 1285
rect 250 1425 360 1450
rect 250 1285 282 1425
rect 328 1285 360 1425
rect 250 1110 360 1285
rect 420 1425 530 1450
rect 420 1285 452 1425
rect 498 1285 530 1425
rect 420 1110 530 1285
rect 590 1425 700 1450
rect 590 1285 622 1425
rect 668 1285 700 1425
rect 590 1110 700 1285
rect 760 1425 860 1450
rect 760 1285 792 1425
rect 838 1285 860 1425
rect 760 1110 860 1285
<< ndiffc >>
rect 142 272 188 318
rect 422 272 468 318
rect 702 272 748 318
<< pdiffc >>
rect 112 1285 158 1425
rect 282 1285 328 1425
rect 452 1285 498 1425
rect 622 1285 668 1425
rect 792 1285 838 1425
<< psubdiff >>
rect 60 118 210 140
rect 60 72 112 118
rect 158 72 210 118
rect 60 50 210 72
rect 290 118 440 140
rect 290 72 342 118
rect 388 72 440 118
rect 290 50 440 72
rect 520 118 670 140
rect 520 72 572 118
rect 618 72 670 118
rect 520 50 670 72
rect 750 118 900 140
rect 750 72 802 118
rect 848 72 900 118
rect 750 50 900 72
<< nsubdiff >>
rect 60 1588 210 1610
rect 60 1542 112 1588
rect 158 1542 210 1588
rect 60 1520 210 1542
rect 290 1588 440 1610
rect 290 1542 342 1588
rect 388 1542 440 1588
rect 290 1520 440 1542
rect 520 1588 670 1610
rect 520 1542 572 1588
rect 618 1542 670 1588
rect 520 1520 670 1542
rect 750 1588 900 1610
rect 750 1542 802 1588
rect 848 1542 900 1588
rect 750 1520 900 1542
<< psubdiffcont >>
rect 112 72 158 118
rect 342 72 388 118
rect 572 72 618 118
rect 802 72 848 118
<< nsubdiffcont >>
rect 112 1542 158 1588
rect 342 1542 388 1588
rect 572 1542 618 1588
rect 802 1542 848 1588
<< polysilicon >>
rect 190 1450 250 1500
rect 360 1450 420 1500
rect 530 1450 590 1500
rect 700 1450 760 1500
rect 190 800 250 1110
rect 360 930 420 1110
rect 300 903 420 930
rect 300 857 347 903
rect 393 857 420 903
rect 300 830 420 857
rect 110 773 250 800
rect 110 727 147 773
rect 193 727 250 773
rect 110 700 250 727
rect 190 490 250 700
rect 360 490 420 830
rect 530 800 590 1110
rect 700 930 760 1110
rect 640 903 760 930
rect 640 857 687 903
rect 733 857 760 903
rect 640 830 760 857
rect 470 773 590 800
rect 470 727 497 773
rect 543 727 590 773
rect 470 700 590 727
rect 530 650 590 700
rect 190 430 280 490
rect 220 380 280 430
rect 330 430 420 490
rect 500 570 590 650
rect 330 380 390 430
rect 500 380 560 570
rect 700 480 760 830
rect 610 420 760 480
rect 610 380 670 420
rect 220 160 280 210
rect 330 160 390 210
rect 500 160 560 210
rect 610 160 670 210
<< polycontact >>
rect 347 857 393 903
rect 147 727 193 773
rect 687 857 733 903
rect 497 727 543 773
<< metal1 >>
rect 0 1588 1070 1660
rect 0 1542 112 1588
rect 158 1542 342 1588
rect 388 1542 572 1588
rect 618 1542 802 1588
rect 848 1542 1070 1588
rect 0 1520 1070 1542
rect 110 1425 160 1450
rect 110 1285 112 1425
rect 158 1285 160 1425
rect 110 1190 160 1285
rect 280 1425 330 1520
rect 280 1285 282 1425
rect 328 1285 330 1425
rect 280 1260 330 1285
rect 450 1425 500 1450
rect 450 1285 452 1425
rect 498 1285 500 1425
rect 620 1425 670 1450
rect 620 1300 622 1425
rect 450 1190 500 1285
rect 600 1285 622 1300
rect 668 1300 670 1425
rect 790 1425 840 1450
rect 668 1296 700 1300
rect 600 1244 624 1285
rect 676 1244 700 1296
rect 600 1240 700 1244
rect 790 1285 792 1425
rect 838 1285 840 1425
rect 790 1190 840 1285
rect 110 1140 840 1190
rect 890 1296 950 1320
rect 890 1244 894 1296
rect 946 1244 950 1296
rect 890 1220 950 1244
rect 890 1040 940 1220
rect 860 1036 960 1040
rect 860 984 884 1036
rect 936 984 960 1036
rect 860 980 960 984
rect 320 906 420 910
rect 320 854 344 906
rect 396 854 420 906
rect 320 850 420 854
rect 660 906 760 910
rect 660 854 684 906
rect 736 854 760 906
rect 660 850 760 854
rect 120 776 220 780
rect 120 724 144 776
rect 196 724 220 776
rect 120 720 220 724
rect 470 776 570 780
rect 470 724 494 776
rect 546 724 570 776
rect 470 720 570 724
rect 880 670 930 980
rect 420 620 930 670
rect 140 318 190 380
rect 140 272 142 318
rect 188 272 190 318
rect 140 140 190 272
rect 420 318 470 620
rect 420 272 422 318
rect 468 272 470 318
rect 420 210 470 272
rect 700 318 750 380
rect 700 272 702 318
rect 748 272 750 318
rect 700 140 750 272
rect 0 118 1070 140
rect 0 72 112 118
rect 158 72 342 118
rect 388 72 572 118
rect 618 72 802 118
rect 848 72 1070 118
rect 0 0 1070 72
<< via1 >>
rect 624 1285 668 1296
rect 668 1285 676 1296
rect 624 1244 676 1285
rect 894 1244 946 1296
rect 884 984 936 1036
rect 344 903 396 906
rect 344 857 347 903
rect 347 857 393 903
rect 393 857 396 903
rect 344 854 396 857
rect 684 903 736 906
rect 684 857 687 903
rect 687 857 733 903
rect 733 857 736 903
rect 684 854 736 857
rect 144 773 196 776
rect 144 727 147 773
rect 147 727 193 773
rect 193 727 196 773
rect 144 724 196 727
rect 494 773 546 776
rect 494 727 497 773
rect 497 727 543 773
rect 543 727 546 773
rect 494 724 546 727
<< metal2 >>
rect 600 1300 700 1310
rect 870 1300 970 1310
rect 600 1296 970 1300
rect 600 1244 624 1296
rect 676 1244 894 1296
rect 946 1244 970 1296
rect 600 1240 970 1244
rect 600 1230 700 1240
rect 870 1230 970 1240
rect 860 1036 960 1050
rect 860 984 884 1036
rect 936 984 960 1036
rect 860 970 960 984
rect 320 906 420 920
rect 320 854 344 906
rect 396 854 420 906
rect 320 840 420 854
rect 660 906 760 920
rect 660 854 684 906
rect 736 854 760 906
rect 660 840 760 854
rect 120 776 220 790
rect 120 724 144 776
rect 196 724 220 776
rect 120 710 220 724
rect 470 776 570 790
rect 470 724 494 776
rect 546 724 570 776
rect 470 710 570 724
<< labels >>
rlabel metal1 s 280 1260 330 1660 4 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 140 0 190 380 4 VSS
port 13 nsew ground bidirectional abutment
rlabel via1 s 894 1244 946 1296 4 Y
port 1 nsew signal output
rlabel via1 s 144 724 196 776 4 A0
port 2 nsew signal input
rlabel via1 s 344 854 396 906 4 A1
port 3 nsew signal input
rlabel via1 s 494 724 546 776 4 B0
port 4 nsew signal input
rlabel via1 s 684 854 736 906 4 B1
port 5 nsew signal input
rlabel metal1 s 0 1520 1070 1660 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 700 0 750 380 1 VSS
port 13 nsew ground bidirectional abutment
rlabel metal1 s 0 0 1070 140 1 VSS
port 13 nsew ground bidirectional abutment
rlabel metal2 s 120 710 220 790 1 A0
port 2 nsew signal input
rlabel metal1 s 120 720 220 780 1 A0
port 2 nsew signal input
rlabel metal2 s 320 840 420 920 1 A1
port 3 nsew signal input
rlabel metal1 s 320 850 420 910 1 A1
port 3 nsew signal input
rlabel metal2 s 470 710 570 790 1 B0
port 4 nsew signal input
rlabel metal1 s 470 720 570 780 1 B0
port 4 nsew signal input
rlabel metal2 s 660 840 760 920 1 B1
port 5 nsew signal input
rlabel metal1 s 660 850 760 910 1 B1
port 5 nsew signal input
rlabel via1 s 884 984 936 1036 1 Y
port 1 nsew signal output
rlabel via1 s 624 1244 676 1296 1 Y
port 1 nsew signal output
rlabel metal2 s 860 970 960 1050 1 Y
port 1 nsew signal output
rlabel metal2 s 600 1230 700 1310 1 Y
port 1 nsew signal output
rlabel metal2 s 600 1240 970 1300 1 Y
port 1 nsew signal output
rlabel metal2 s 870 1230 970 1310 1 Y
port 1 nsew signal output
rlabel metal1 s 620 1240 670 1450 1 Y
port 1 nsew signal output
rlabel metal1 s 600 1240 700 1300 1 Y
port 1 nsew signal output
rlabel metal1 s 420 210 470 670 1 Y
port 1 nsew signal output
rlabel metal1 s 420 620 930 670 1 Y
port 1 nsew signal output
rlabel metal1 s 880 620 930 1040 1 Y
port 1 nsew signal output
rlabel metal1 s 890 980 940 1320 1 Y
port 1 nsew signal output
rlabel metal1 s 890 1220 950 1320 1 Y
port 1 nsew signal output
rlabel metal1 s 860 980 960 1040 1 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1070 1660
string GDS_END 48216
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_gp12t3v3/gds/gf180mcu_osu_sc_gp12t3v3.gds
string GDS_START 41414
string LEFclass CORE
string LEFsite gf180mcu_osu_sc_gp12t3v3
string LEFsymmetry X Y
<< end >>
