VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__fillnc
  CLASS PAD SPACER ;
  FOREIGN gf180mcu_fd_io__fillnc ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.100 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 0.100 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 0.100 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 0.100 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 0.100 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 0.100 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 0.100 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 0.100 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 0.100 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 0.100 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 0.100 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 0.100 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 0.100 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 0.100 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 0.100 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 0.100 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 0.100 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 0.100 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 0.100 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 0.100 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 0.100 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 0.100 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 0.100 85.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 0.100 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 0.100 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 0.100 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 0.100 253.000 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 0.260 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 246.000 0.100 325.000 ;
  END
END gf180mcu_fd_io__fillnc
END LIBRARY

